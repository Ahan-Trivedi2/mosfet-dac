magic
tech sky130A
<< checkpaint >>
rect 19714 15016 27656 15286
rect 19694 14826 27656 15016
rect 19444 14786 27656 14826
rect 19444 14046 27806 14786
rect 19444 13956 28116 14046
rect 19444 13306 28506 13956
rect 14774 11306 28506 13306
rect -1996 6876 5936 6906
rect -1996 -2006 11136 6876
rect 3204 -2076 11136 -2006
rect 14774 3536 32736 11306
rect 14774 2376 33826 3536
rect 14774 -574 34246 2376
rect 14774 -4944 35216 -574
rect 7994 -5636 35216 -4944
rect 7994 -6406 34326 -5636
rect 7994 -6516 30526 -6406
rect 7994 -8646 27656 -6516
rect 7994 -10006 16646 -8646
rect 8544 -10876 14676 -10006
rect 19594 -10746 27656 -8646
rect 8544 -12256 13276 -10876
rect 8544 -12666 12766 -12256
rect 19714 -12306 27656 -10746
<< nwell >>
rect 18290 -1380 18310 -1140
rect 18830 -1380 18850 -1140
rect 19370 -1380 19390 -1140
rect 19910 -1380 19930 -1140
<< locali >>
rect 17350 -1050 17400 -1040
rect 17350 -1130 17360 -1050
rect 17390 -1130 17400 -1050
rect 17350 -1140 17400 -1130
rect 17520 -1050 17570 -1040
rect 17520 -1130 17530 -1050
rect 17560 -1130 17570 -1050
rect 17520 -1640 17570 -1130
rect 17890 -1050 17940 -1040
rect 17890 -1130 17900 -1050
rect 17930 -1130 17940 -1050
rect 17890 -1140 17940 -1130
rect 18060 -1050 18110 -1040
rect 18060 -1130 18070 -1050
rect 18100 -1130 18110 -1050
rect 18060 -1640 18110 -1130
rect 18430 -1050 18480 -1040
rect 18430 -1130 18440 -1050
rect 18470 -1130 18480 -1050
rect 18430 -1140 18480 -1130
rect 18600 -1050 18650 -1040
rect 18600 -1130 18610 -1050
rect 18640 -1130 18650 -1050
rect 18600 -1640 18650 -1130
rect 18970 -1050 19020 -1040
rect 18970 -1130 18980 -1050
rect 19010 -1130 19020 -1050
rect 18970 -1140 19020 -1130
rect 19140 -1050 19190 -1040
rect 19140 -1130 19150 -1050
rect 19180 -1130 19190 -1050
rect 19140 -1640 19190 -1130
rect 19510 -1050 19560 -1040
rect 19510 -1130 19520 -1050
rect 19550 -1130 19560 -1050
rect 19510 -1140 19560 -1130
rect 19680 -1050 19730 -1040
rect 19680 -1130 19690 -1050
rect 19720 -1130 19730 -1050
rect 19680 -1640 19730 -1130
rect 20050 -1050 20100 -1040
rect 20050 -1130 20060 -1050
rect 20090 -1130 20100 -1050
rect 20050 -1140 20100 -1130
rect 20220 -1050 20270 -1040
rect 20220 -1130 20230 -1050
rect 20260 -1130 20270 -1050
rect 20220 -1640 20270 -1130
rect 17520 -1680 17770 -1640
rect 18060 -1680 18310 -1640
rect 18600 -1680 18850 -1640
rect 19140 -1680 19390 -1640
rect 19680 -1680 19930 -1640
rect 20220 -1680 20470 -1640
<< viali >>
rect 17360 -1130 17390 -1050
rect 17530 -1130 17560 -1050
rect 17900 -1130 17930 -1050
rect 18070 -1130 18100 -1050
rect 18440 -1130 18470 -1050
rect 18610 -1130 18640 -1050
rect 18980 -1130 19010 -1050
rect 19150 -1130 19180 -1050
rect 19520 -1130 19550 -1050
rect 19690 -1130 19720 -1050
rect 20060 -1130 20090 -1050
rect 20230 -1130 20260 -1050
<< metal1 >>
rect 17350 -1045 17400 -1040
rect 17350 -1135 17355 -1045
rect 17395 -1135 17400 -1045
rect 17350 -1140 17400 -1135
rect 17520 -1045 17570 -1040
rect 17520 -1135 17525 -1045
rect 17565 -1135 17570 -1045
rect 17520 -1140 17570 -1135
rect 17890 -1045 17940 -1040
rect 17890 -1135 17895 -1045
rect 17935 -1135 17940 -1045
rect 17890 -1140 17940 -1135
rect 18060 -1045 18110 -1040
rect 18060 -1135 18065 -1045
rect 18105 -1135 18110 -1045
rect 18060 -1140 18110 -1135
rect 18430 -1045 18480 -1040
rect 18430 -1135 18435 -1045
rect 18475 -1135 18480 -1045
rect 18430 -1140 18480 -1135
rect 18600 -1045 18650 -1040
rect 18600 -1135 18605 -1045
rect 18645 -1135 18650 -1045
rect 18600 -1140 18650 -1135
rect 18970 -1045 19020 -1040
rect 18970 -1135 18975 -1045
rect 19015 -1135 19020 -1045
rect 18970 -1140 19020 -1135
rect 19140 -1045 19190 -1040
rect 19140 -1135 19145 -1045
rect 19185 -1135 19190 -1045
rect 19140 -1140 19190 -1135
rect 19510 -1045 19560 -1040
rect 19510 -1135 19515 -1045
rect 19555 -1135 19560 -1045
rect 19510 -1140 19560 -1135
rect 19680 -1045 19730 -1040
rect 19680 -1135 19685 -1045
rect 19725 -1135 19730 -1045
rect 19680 -1140 19730 -1135
rect 20050 -1045 20100 -1040
rect 20050 -1135 20055 -1045
rect 20095 -1135 20100 -1045
rect 20050 -1140 20100 -1135
rect 20220 -1045 20270 -1040
rect 20220 -1135 20225 -1045
rect 20265 -1135 20270 -1045
rect 20220 -1140 20270 -1135
<< via1 >>
rect 17355 -1050 17395 -1045
rect 17355 -1130 17360 -1050
rect 17360 -1130 17390 -1050
rect 17390 -1130 17395 -1050
rect 17355 -1135 17395 -1130
rect 17525 -1050 17565 -1045
rect 17525 -1130 17530 -1050
rect 17530 -1130 17560 -1050
rect 17560 -1130 17565 -1050
rect 17525 -1135 17565 -1130
rect 17895 -1050 17935 -1045
rect 17895 -1130 17900 -1050
rect 17900 -1130 17930 -1050
rect 17930 -1130 17935 -1050
rect 17895 -1135 17935 -1130
rect 18065 -1050 18105 -1045
rect 18065 -1130 18070 -1050
rect 18070 -1130 18100 -1050
rect 18100 -1130 18105 -1050
rect 18065 -1135 18105 -1130
rect 18435 -1050 18475 -1045
rect 18435 -1130 18440 -1050
rect 18440 -1130 18470 -1050
rect 18470 -1130 18475 -1050
rect 18435 -1135 18475 -1130
rect 18605 -1050 18645 -1045
rect 18605 -1130 18610 -1050
rect 18610 -1130 18640 -1050
rect 18640 -1130 18645 -1050
rect 18605 -1135 18645 -1130
rect 18975 -1050 19015 -1045
rect 18975 -1130 18980 -1050
rect 18980 -1130 19010 -1050
rect 19010 -1130 19015 -1050
rect 18975 -1135 19015 -1130
rect 19145 -1050 19185 -1045
rect 19145 -1130 19150 -1050
rect 19150 -1130 19180 -1050
rect 19180 -1130 19185 -1050
rect 19145 -1135 19185 -1130
rect 19515 -1050 19555 -1045
rect 19515 -1130 19520 -1050
rect 19520 -1130 19550 -1050
rect 19550 -1130 19555 -1050
rect 19515 -1135 19555 -1130
rect 19685 -1050 19725 -1045
rect 19685 -1130 19690 -1050
rect 19690 -1130 19720 -1050
rect 19720 -1130 19725 -1050
rect 19685 -1135 19725 -1130
rect 20055 -1050 20095 -1045
rect 20055 -1130 20060 -1050
rect 20060 -1130 20090 -1050
rect 20090 -1130 20095 -1050
rect 20055 -1135 20095 -1130
rect 20225 -1050 20265 -1045
rect 20225 -1130 20230 -1050
rect 20230 -1130 20260 -1050
rect 20260 -1130 20265 -1050
rect 20225 -1135 20265 -1130
<< metal2 >>
rect 17350 -1045 17400 -1040
rect 17350 -1135 17355 -1045
rect 17395 -1135 17400 -1045
rect 17350 -1140 17400 -1135
rect 17520 -1045 17570 -1040
rect 17520 -1135 17525 -1045
rect 17565 -1135 17570 -1045
rect 17520 -1140 17570 -1135
rect 17890 -1045 17940 -1040
rect 17890 -1135 17895 -1045
rect 17935 -1135 17940 -1045
rect 17890 -1140 17940 -1135
rect 18060 -1045 18110 -1040
rect 18060 -1135 18065 -1045
rect 18105 -1135 18110 -1045
rect 18060 -1140 18110 -1135
rect 18430 -1045 18480 -1040
rect 18430 -1135 18435 -1045
rect 18475 -1135 18480 -1045
rect 18430 -1140 18480 -1135
rect 18600 -1045 18650 -1040
rect 18600 -1135 18605 -1045
rect 18645 -1135 18650 -1045
rect 18600 -1140 18650 -1135
rect 18970 -1045 19020 -1040
rect 18970 -1135 18975 -1045
rect 19015 -1135 19020 -1045
rect 18970 -1140 19020 -1135
rect 19140 -1045 19190 -1040
rect 19140 -1135 19145 -1045
rect 19185 -1135 19190 -1045
rect 19140 -1140 19190 -1135
rect 19510 -1045 19560 -1040
rect 19510 -1135 19515 -1045
rect 19555 -1135 19560 -1045
rect 19510 -1140 19560 -1135
rect 19680 -1045 19730 -1040
rect 19680 -1135 19685 -1045
rect 19725 -1135 19730 -1045
rect 19680 -1140 19730 -1135
rect 20050 -1045 20100 -1040
rect 20050 -1135 20055 -1045
rect 20095 -1135 20100 -1045
rect 20050 -1140 20100 -1135
rect 20220 -1045 20270 -1040
rect 20220 -1135 20225 -1045
rect 20265 -1135 20270 -1045
rect 20220 -1140 20270 -1135
<< via2 >>
rect 17355 -1135 17395 -1045
rect 17525 -1135 17565 -1045
rect 17895 -1135 17935 -1045
rect 18065 -1135 18105 -1045
rect 18435 -1135 18475 -1045
rect 18605 -1135 18645 -1045
rect 18975 -1135 19015 -1045
rect 19145 -1135 19185 -1045
rect 19515 -1135 19555 -1045
rect 19685 -1135 19725 -1045
rect 20055 -1135 20095 -1045
rect 20225 -1135 20265 -1045
<< metal3 >>
rect 17350 -1045 17400 -1040
rect 17350 -1135 17355 -1045
rect 17395 -1135 17400 -1045
rect 17350 -1140 17400 -1135
rect 17520 -1045 17570 -1040
rect 17520 -1135 17525 -1045
rect 17565 -1135 17570 -1045
rect 17520 -1140 17570 -1135
rect 17890 -1045 17940 -1040
rect 17890 -1135 17895 -1045
rect 17935 -1135 17940 -1045
rect 17890 -1140 17940 -1135
rect 18060 -1045 18110 -1040
rect 18060 -1135 18065 -1045
rect 18105 -1135 18110 -1045
rect 18060 -1140 18110 -1135
rect 18430 -1045 18480 -1040
rect 18430 -1135 18435 -1045
rect 18475 -1135 18480 -1045
rect 18430 -1140 18480 -1135
rect 18600 -1045 18650 -1040
rect 18600 -1135 18605 -1045
rect 18645 -1135 18650 -1045
rect 18600 -1140 18650 -1135
rect 18970 -1045 19020 -1040
rect 18970 -1135 18975 -1045
rect 19015 -1135 19020 -1045
rect 18970 -1140 19020 -1135
rect 19140 -1045 19190 -1040
rect 19140 -1135 19145 -1045
rect 19185 -1135 19190 -1045
rect 19140 -1140 19190 -1135
rect 19510 -1045 19560 -1040
rect 19510 -1135 19515 -1045
rect 19555 -1135 19560 -1045
rect 19510 -1140 19560 -1135
rect 19680 -1045 19730 -1040
rect 19680 -1135 19685 -1045
rect 19725 -1135 19730 -1045
rect 19680 -1140 19730 -1135
rect 20050 -1045 20100 -1040
rect 20050 -1135 20055 -1045
rect 20095 -1135 20100 -1045
rect 20050 -1140 20100 -1135
rect 20220 -1045 20270 -1040
rect 20220 -1135 20225 -1045
rect 20265 -1135 20270 -1045
rect 20220 -1140 20270 -1135
use bbg  bbg_0
timestamp 1762117721
transform 1 0 21910 0 1 -2470
box -220 -560 1820 210
use ccm  ccm_0
timestamp 1762061669
transform 0 1 23990 -1 0 -660
box -1810 -10 2910 1120
use dac  dac_0
timestamp 1762117972
transform 1 0 17190 0 1 7535
box -450 -8595 4340 3805
use fvf  fvf_0
timestamp 1762123188
transform 0 1 23360 -1 0 1005
box -150 -510 3125 510
use fvf  fvf_1
timestamp 1762123188
transform 0 1 22210 -1 0 1005
box -150 -510 3125 510
use inv  inv_0
timestamp 1762145583
transform 1 0 17300 0 1 -1630
box -90 -50 200 490
use inv  inv_1
timestamp 1762145583
transform 1 0 17840 0 1 -1630
box -90 -50 200 490
use inv  inv_2
timestamp 1762145583
transform 1 0 18380 0 1 -1630
box -90 -50 200 490
use inv  inv_3
timestamp 1762145583
transform 1 0 18920 0 1 -1630
box -90 -50 200 490
use inv  inv_4
timestamp 1762145583
transform 1 0 19460 0 1 -1630
box -90 -50 200 490
use inv  inv_5
timestamp 1762145583
transform 1 0 20000 0 1 -1630
box -90 -50 200 490
use inv  inv_6
timestamp 1762145583
transform 1 0 20540 0 1 -1630
box -90 -50 200 490
use ncbc  ncbc_0
timestamp 1762057603
transform 1 0 22010 0 1 450
box -310 810 3690 5830
use pcbc  pcbc_0
timestamp 1762057942
transform 1 0 17560 0 1 3680
box 4150 2710 8150 7690
<< end >>
