magic
tech sky130A
timestamp 1762205191
<< nwell >>
rect 2030 11130 2500 11380
rect 3260 11130 3730 11380
rect 2350 7090 2490 7370
<< nmos >>
rect 2580 11270 2680 11370
rect 2720 11270 2820 11370
rect 2940 11270 3040 11370
rect 3080 11270 3180 11370
rect 2580 11140 2680 11240
rect 2720 11140 2820 11240
rect 2940 11140 3040 11240
rect 3080 11140 3180 11240
<< pmos >>
rect 2140 11290 2440 11345
rect 3320 11290 3620 11345
rect 2140 11160 2440 11215
rect 3320 11160 3620 11215
rect 2370 7200 2470 7300
<< ndiff >>
rect 2540 11340 2580 11370
rect 2540 11300 2550 11340
rect 2570 11300 2580 11340
rect 2540 11270 2580 11300
rect 2680 11340 2720 11370
rect 2680 11300 2690 11340
rect 2710 11300 2720 11340
rect 2680 11270 2720 11300
rect 2820 11340 2860 11370
rect 2900 11340 2940 11370
rect 2820 11300 2830 11340
rect 2850 11300 2860 11340
rect 2900 11300 2910 11340
rect 2930 11300 2940 11340
rect 2820 11270 2860 11300
rect 2900 11270 2940 11300
rect 3040 11340 3080 11370
rect 3040 11300 3050 11340
rect 3070 11300 3080 11340
rect 3040 11270 3080 11300
rect 3180 11340 3220 11370
rect 3180 11300 3190 11340
rect 3210 11300 3220 11340
rect 3180 11270 3220 11300
rect 2540 11210 2580 11240
rect 2540 11170 2550 11210
rect 2570 11170 2580 11210
rect 2540 11140 2580 11170
rect 2680 11210 2720 11240
rect 2680 11170 2690 11210
rect 2710 11170 2720 11210
rect 2680 11140 2720 11170
rect 2820 11210 2860 11240
rect 2900 11210 2940 11240
rect 2820 11170 2830 11210
rect 2850 11170 2860 11210
rect 2900 11170 2910 11210
rect 2930 11170 2940 11210
rect 2820 11140 2860 11170
rect 2900 11140 2940 11170
rect 3040 11210 3080 11240
rect 3040 11170 3050 11210
rect 3070 11170 3080 11210
rect 3040 11140 3080 11170
rect 3180 11210 3220 11240
rect 3180 11170 3190 11210
rect 3210 11170 3220 11210
rect 3180 11140 3220 11170
<< pdiff >>
rect 2100 11340 2140 11345
rect 2100 11300 2110 11340
rect 2130 11300 2140 11340
rect 2100 11290 2140 11300
rect 2440 11340 2480 11345
rect 2440 11300 2450 11340
rect 2470 11300 2480 11340
rect 2440 11290 2480 11300
rect 3280 11340 3320 11345
rect 3280 11300 3290 11340
rect 3310 11300 3320 11340
rect 3280 11290 3320 11300
rect 3620 11340 3660 11345
rect 3620 11300 3630 11340
rect 3650 11300 3660 11340
rect 3620 11290 3660 11300
rect 2100 11210 2140 11215
rect 2100 11170 2110 11210
rect 2130 11170 2140 11210
rect 2100 11160 2140 11170
rect 2440 11210 2480 11215
rect 2440 11170 2450 11210
rect 2470 11170 2480 11210
rect 2440 11160 2480 11170
rect 3280 11210 3320 11215
rect 3280 11170 3290 11210
rect 3310 11170 3320 11210
rect 3280 11160 3320 11170
rect 3620 11210 3660 11215
rect 3620 11170 3630 11210
rect 3650 11170 3660 11210
rect 3620 11160 3660 11170
rect 2370 7340 2470 7350
rect 2370 7310 2390 7340
rect 2450 7310 2470 7340
rect 2370 7300 2470 7310
rect 2370 7190 2470 7200
rect 2370 7160 2390 7190
rect 2450 7160 2470 7190
rect 2370 7150 2470 7160
<< ndiffc >>
rect 2550 11300 2570 11340
rect 2690 11300 2710 11340
rect 2830 11300 2850 11340
rect 2910 11300 2930 11340
rect 3050 11300 3070 11340
rect 3190 11300 3210 11340
rect 2550 11170 2570 11210
rect 2690 11170 2710 11210
rect 2830 11170 2850 11210
rect 2910 11170 2930 11210
rect 3050 11170 3070 11210
rect 3190 11170 3210 11210
<< pdiffc >>
rect 2110 11300 2130 11340
rect 2450 11300 2470 11340
rect 3290 11300 3310 11340
rect 3630 11300 3650 11340
rect 2110 11170 2130 11210
rect 2450 11170 2470 11210
rect 3290 11170 3310 11210
rect 3630 11170 3650 11210
rect 2390 7310 2450 7340
rect 2390 7160 2450 7190
<< psubdiff >>
rect 2860 11340 2900 11370
rect 2860 11300 2870 11340
rect 2890 11300 2900 11340
rect 2860 11270 2900 11300
rect 2860 11210 2900 11240
rect 2860 11170 2870 11210
rect 2890 11170 2900 11210
rect 2860 11140 2900 11170
<< nsubdiff >>
rect 2050 11345 2080 11360
rect 2050 11340 2100 11345
rect 2050 11300 2070 11340
rect 2090 11300 2100 11340
rect 2050 11290 2100 11300
rect 2050 11280 2080 11290
rect 2050 11215 2080 11230
rect 3680 11345 3710 11360
rect 3660 11340 3710 11345
rect 3660 11300 3670 11340
rect 3690 11300 3710 11340
rect 3660 11290 3710 11300
rect 2050 11210 2100 11215
rect 2050 11170 2070 11210
rect 2090 11170 2100 11210
rect 2050 11160 2100 11170
rect 2050 11150 2080 11160
rect 3680 11280 3710 11290
rect 3680 11215 3710 11230
rect 3660 11210 3710 11215
rect 3660 11170 3670 11210
rect 3690 11170 3710 11210
rect 3660 11160 3710 11170
rect 3680 11150 3710 11160
rect 2370 7140 2470 7150
rect 2370 7110 2390 7140
rect 2450 7110 2470 7140
<< psubdiffcont >>
rect 2870 11300 2890 11340
rect 2870 11170 2890 11210
<< nsubdiffcont >>
rect 2070 11300 2090 11340
rect 3670 11300 3690 11340
rect 2070 11170 2090 11210
rect 3670 11170 3690 11210
rect 2390 7110 2450 7140
<< poly >>
rect 2580 11370 2680 11390
rect 2720 11370 2820 11390
rect 2940 11370 3040 11390
rect 3080 11370 3180 11390
rect 2140 11345 2440 11370
rect 2140 11215 2440 11290
rect 3320 11345 3620 11370
rect 2580 11240 2680 11270
rect 2720 11240 2820 11270
rect 2940 11240 3040 11270
rect 3080 11240 3180 11270
rect 2140 11140 2440 11160
rect 3320 11215 3620 11290
rect 3320 11140 3620 11160
rect 2140 11130 2180 11140
rect 2140 11110 2150 11130
rect 2170 11110 2180 11130
rect 2140 11100 2180 11110
rect 2580 11120 2680 11140
rect 2720 11120 2820 11140
rect 2940 11120 3040 11140
rect 3080 11120 3180 11140
rect 2580 11100 2590 11120
rect 2610 11100 2620 11120
rect 2580 11090 2620 11100
rect 2720 11100 2730 11120
rect 2750 11100 2760 11120
rect 2720 11090 2760 11100
rect 3000 11100 3010 11120
rect 3030 11100 3040 11120
rect 3000 11090 3040 11100
rect 3140 11100 3150 11120
rect 3170 11100 3180 11120
rect 3580 11130 3620 11140
rect 3580 11110 3590 11130
rect 3610 11110 3620 11130
rect 3580 11100 3620 11110
rect 3140 11090 3180 11100
rect 2280 7270 2370 7300
rect 2280 7230 2300 7270
rect 2340 7230 2370 7270
rect 2280 7200 2370 7230
rect 2470 7200 2490 7300
rect 9720 55 9765 70
rect 9725 35 9735 55
rect 9755 35 9765 55
rect 9725 25 9765 35
<< polycont >>
rect 2150 11110 2170 11130
rect 2590 11100 2610 11120
rect 2730 11100 2750 11120
rect 3010 11100 3030 11120
rect 3150 11100 3170 11120
rect 3590 11110 3610 11130
rect 2300 7230 2340 7270
rect 9735 35 9755 55
<< locali >>
rect 1700 7400 1750 13590
rect 2100 11450 3660 11470
rect 2050 11345 2080 11360
rect 2100 11345 2140 11450
rect 2540 11410 3220 11430
rect 2540 11350 2580 11410
rect 2480 11345 2580 11350
rect 2050 11340 2140 11345
rect 2050 11300 2070 11340
rect 2090 11300 2110 11340
rect 2130 11300 2140 11340
rect 2050 11290 2140 11300
rect 2440 11340 2580 11345
rect 2440 11300 2450 11340
rect 2470 11300 2550 11340
rect 2570 11300 2580 11340
rect 2440 11290 2580 11300
rect 2050 11280 2080 11290
rect 2050 11215 2080 11230
rect 2100 11215 2140 11290
rect 2540 11220 2580 11290
rect 2480 11215 2580 11220
rect 2050 11210 2140 11215
rect 2050 11170 2070 11210
rect 2090 11170 2110 11210
rect 2130 11170 2140 11210
rect 2050 11160 2140 11170
rect 2440 11210 2580 11215
rect 2440 11170 2450 11210
rect 2470 11170 2550 11210
rect 2570 11170 2580 11210
rect 2440 11160 2580 11170
rect 2050 11150 2080 11160
rect 2140 11130 2180 11140
rect 2140 11110 2150 11130
rect 2170 11110 2180 11130
rect 2140 11100 2180 11110
rect 2540 11130 2580 11160
rect 2680 11370 3080 11390
rect 2680 11340 2720 11370
rect 2680 11300 2690 11340
rect 2710 11300 2720 11340
rect 2680 11210 2720 11300
rect 2680 11170 2690 11210
rect 2710 11170 2720 11210
rect 2680 11130 2720 11170
rect 2820 11340 2940 11350
rect 2820 11300 2830 11340
rect 2850 11300 2870 11340
rect 2890 11300 2910 11340
rect 2930 11300 2940 11340
rect 2820 11210 2940 11300
rect 2820 11170 2830 11210
rect 2850 11170 2870 11210
rect 2890 11170 2910 11210
rect 2930 11170 2940 11210
rect 2540 11120 2620 11130
rect 2540 11100 2590 11120
rect 2610 11100 2620 11120
rect 2540 11090 2620 11100
rect 2680 11120 2760 11130
rect 2680 11100 2730 11120
rect 2750 11100 2760 11120
rect 2680 11090 2760 11100
rect 2820 11090 2940 11170
rect 3040 11340 3080 11370
rect 3040 11300 3050 11340
rect 3070 11300 3080 11340
rect 3040 11210 3080 11300
rect 3040 11170 3050 11210
rect 3070 11170 3080 11210
rect 3040 11130 3080 11170
rect 3180 11350 3220 11410
rect 3180 11345 3280 11350
rect 3620 11345 3660 11450
rect 3680 11345 3710 11360
rect 3180 11340 3320 11345
rect 3180 11300 3190 11340
rect 3210 11300 3290 11340
rect 3310 11300 3320 11340
rect 3180 11290 3320 11300
rect 3620 11340 3710 11345
rect 3620 11300 3630 11340
rect 3650 11300 3670 11340
rect 3690 11300 3710 11340
rect 3620 11290 3710 11300
rect 3180 11220 3220 11290
rect 3180 11215 3280 11220
rect 3620 11215 3660 11290
rect 3680 11280 3710 11290
rect 3680 11215 3710 11230
rect 3180 11210 3320 11215
rect 3180 11170 3190 11210
rect 3210 11170 3290 11210
rect 3310 11170 3320 11210
rect 3180 11160 3320 11170
rect 3620 11210 3710 11215
rect 3620 11170 3630 11210
rect 3650 11170 3670 11210
rect 3690 11170 3710 11210
rect 3620 11160 3710 11170
rect 3180 11130 3220 11160
rect 3000 11120 3080 11130
rect 3000 11100 3010 11120
rect 3030 11100 3080 11120
rect 3000 11090 3080 11100
rect 3140 11120 3220 11130
rect 3140 11100 3150 11120
rect 3170 11100 3220 11120
rect 3580 11130 3620 11140
rect 3580 11110 3590 11130
rect 3610 11110 3620 11130
rect 3580 11100 3620 11110
rect 3140 11090 3220 11100
rect 2820 10830 2860 11090
rect 3660 11040 3710 11160
rect 2780 10780 2860 10830
rect 3620 10980 3710 11040
rect 2780 10670 2820 10780
rect 2770 10660 2820 10670
rect 2770 10640 2780 10660
rect 2810 10640 2820 10660
rect 2770 10630 2820 10640
rect 3620 10610 3660 10980
rect 2560 10550 3660 10610
rect 1700 7350 2460 7400
rect 2380 7340 2460 7350
rect 2380 7310 2390 7340
rect 2450 7310 2460 7340
rect 2380 7300 2460 7310
rect 2280 7270 2360 7300
rect 2280 7230 2300 7270
rect 2340 7230 2360 7270
rect 2280 7200 2360 7230
rect 2560 7200 2630 10550
rect 2770 10510 2810 10520
rect 2770 10480 2780 10510
rect 2800 10480 2810 10510
rect 2770 7750 2810 10480
rect 6865 7905 6945 7910
rect 6865 7885 6870 7905
rect 6940 7885 6945 7905
rect 6865 7875 6945 7885
rect 2770 7710 2780 7750
rect 2800 7710 2810 7750
rect 2770 7690 2810 7710
rect 2380 7190 2620 7200
rect 2380 7160 2390 7190
rect 2450 7160 2620 7190
rect 2380 7150 2620 7160
rect 2370 7140 2470 7150
rect 2370 7110 2390 7140
rect 2450 7110 2470 7140
rect 6800 5380 7150 5420
rect 6800 5315 6915 5325
rect 6800 5295 6810 5315
rect 6880 5295 6915 5315
rect 6800 5285 6915 5295
rect 1310 1480 1350 4780
rect 1300 1460 1350 1480
rect 1300 1430 1310 1460
rect 1340 1430 1350 1460
rect 1300 1420 1350 1430
rect 7100 1370 7150 5380
rect 8400 3440 8430 3450
rect 8500 3440 8530 3450
rect 8400 3435 8530 3440
rect 8400 3410 8405 3435
rect 8425 3410 8505 3435
rect 8525 3410 8530 3435
rect 8400 3400 8530 3410
rect 8400 3340 8430 3350
rect 8500 3340 8530 3350
rect 8400 3335 8530 3340
rect 8400 3310 8405 3335
rect 8425 3310 8505 3335
rect 8525 3310 8530 3335
rect 8400 3300 8530 3310
rect 7100 1320 9230 1370
rect 7110 1230 9120 1270
rect -3040 680 -3020 1020
rect -2260 880 -2240 1010
rect -2300 850 -2240 880
rect -2300 830 -2270 850
rect -2080 830 -2060 1020
rect -1710 880 -1690 1030
rect -1540 880 -1520 1010
rect -1170 930 -1150 1000
rect -1000 930 -980 1000
rect -630 930 -610 1000
rect -460 930 -440 1000
rect -100 980 -80 1000
rect -1230 900 -1150 930
rect -1030 900 -980 930
rect -780 900 -610 930
rect -580 900 -440 930
rect -250 950 -80 980
rect -1230 880 -1200 900
rect -1030 880 -1000 900
rect -780 880 -750 900
rect -580 880 -550 900
rect -250 880 -220 950
rect 80 930 100 990
rect -1850 850 -1690 880
rect -1600 850 -1520 880
rect -1400 850 -1200 880
rect -1180 850 -1000 880
rect -980 850 -750 880
rect -730 850 -550 880
rect -530 850 -220 880
rect -200 900 100 930
rect 450 920 470 980
rect -1850 830 -1820 850
rect -1600 830 -1570 850
rect -1400 830 -1370 850
rect -1180 830 -1150 850
rect -980 830 -950 850
rect -730 830 -700 850
rect -530 830 -500 850
rect -200 830 -170 900
rect 170 890 470 920
rect 170 880 210 890
rect -2450 800 -2270 830
rect -2250 800 -2060 830
rect -2000 800 -1820 830
rect -1800 800 -1570 830
rect -1550 800 -1370 830
rect -1350 800 -1150 830
rect -1130 800 -950 830
rect -930 800 -700 830
rect -680 800 -500 830
rect -480 800 -170 830
rect -150 850 210 880
rect 620 870 640 990
rect -2450 780 -2420 800
rect -2250 780 -2220 800
rect -2000 780 -1970 800
rect -1800 780 -1770 800
rect -1550 780 -1520 800
rect -1350 780 -1320 800
rect -1130 780 -1100 800
rect -930 780 -900 800
rect -680 780 -650 800
rect -480 780 -450 800
rect -150 780 -120 850
rect 230 840 640 870
rect 230 830 270 840
rect -2650 750 -2420 780
rect -2400 750 -2220 780
rect -2200 750 -1970 780
rect -1950 750 -1770 780
rect -1750 750 -1520 780
rect -1500 750 -1320 780
rect -1300 750 -1100 780
rect -1080 750 -900 780
rect -880 750 -650 780
rect -630 750 -450 780
rect -430 750 -120 780
rect -100 800 270 830
rect 1140 820 1160 990
rect -2650 730 -2620 750
rect -2400 730 -2370 750
rect -2200 730 -2170 750
rect -1950 730 -1920 750
rect -1750 730 -1720 750
rect -1500 730 -1470 750
rect -1300 730 -1270 750
rect -1080 730 -1050 750
rect -880 730 -850 750
rect -630 730 -600 750
rect -430 730 -400 750
rect -100 730 -70 800
rect 290 790 1160 820
rect 2040 830 2080 840
rect 290 780 330 790
rect -2800 700 -2620 730
rect -2600 700 -2370 730
rect -2350 700 -2170 730
rect -2150 700 -1920 730
rect -1900 700 -1720 730
rect -1700 700 -1470 730
rect -1450 700 -1270 730
rect -1250 700 -1050 730
rect -1030 700 -850 730
rect -830 700 -600 730
rect -580 700 -400 730
rect -380 700 -70 730
rect -50 750 330 780
rect 2040 760 2050 830
rect 2070 760 2080 830
rect 2040 750 2080 760
rect 2195 830 2235 840
rect 2195 760 2205 830
rect 2225 760 2235 830
rect -2800 680 -2770 700
rect -2600 680 -2570 700
rect -2350 680 -2320 700
rect -2150 680 -2120 700
rect -1900 680 -1870 700
rect -1700 680 -1670 700
rect -1450 680 -1420 700
rect -1250 680 -1220 700
rect -1030 680 -1000 700
rect -830 680 -800 700
rect -580 680 -550 700
rect -380 680 -350 700
rect -50 680 -20 750
rect -3170 650 -3020 680
rect -2970 650 -2770 680
rect -2750 650 -2570 680
rect -2550 650 -2320 680
rect -2300 650 -2120 680
rect -2100 650 -1870 680
rect -1850 650 -1670 680
rect -1650 650 -1420 680
rect -1400 650 -1220 680
rect -1200 650 -1000 680
rect -980 650 -800 680
rect -780 650 -550 680
rect -530 650 -350 680
rect -330 650 -20 680
rect -3170 150 -3130 650
rect -2750 150 -2710 650
rect -2300 150 -2260 650
rect -1850 150 -1810 650
rect -1400 150 -1360 650
rect -980 150 -940 650
rect -530 150 -490 650
rect -330 640 -290 650
rect -3170 110 -3090 150
rect -2750 110 -2670 150
rect -2300 110 -2220 150
rect -1850 110 -1770 150
rect -1400 110 -1320 150
rect -980 110 -900 150
rect -530 110 -450 150
rect 2195 40 2235 760
rect 7110 160 7150 1230
rect 9080 1130 9120 1230
rect 9180 1260 9230 1320
rect 9180 1230 9190 1260
rect 9220 1230 9230 1260
rect 9180 1210 9230 1230
rect 10650 1080 10720 1820
rect 10500 1040 10720 1080
rect 6800 120 7150 160
rect 9725 60 9765 70
rect 2040 20 2235 40
rect 9725 30 9730 60
rect 9760 30 9765 60
rect 9725 25 9765 30
<< viali >>
rect 2550 11300 2570 11340
rect 2150 11110 2170 11130
rect 3590 11110 3610 11130
rect 2780 10640 2810 10660
rect 2390 7310 2450 7340
rect 2300 7230 2340 7270
rect 2780 10480 2800 10510
rect 6870 7885 6940 7905
rect 2780 7710 2800 7750
rect 2390 7160 2450 7190
rect 2870 5295 2940 5315
rect 6810 5295 6880 5315
rect 1310 1430 1340 1460
rect 8405 3410 8425 3435
rect 8505 3410 8525 3435
rect 8405 3310 8425 3335
rect 8505 3310 8525 3335
rect 2050 760 2070 830
rect 2205 760 2225 830
rect -3090 520 -3070 540
rect -3090 250 -3070 270
rect -2670 520 -2650 540
rect -2670 250 -2650 270
rect -2220 520 -2200 540
rect -2220 250 -2200 270
rect -1770 520 -1750 540
rect -1770 250 -1750 270
rect -1320 520 -1300 540
rect -1320 250 -1300 270
rect -900 520 -880 540
rect -900 250 -880 270
rect -450 520 -430 540
rect -450 250 -430 270
rect 9190 1230 9220 1260
rect 7510 970 7540 1000
rect 9800 380 9830 410
rect 2840 25 2910 45
rect 9190 30 9220 60
rect 9730 55 9760 60
rect 9730 35 9735 55
rect 9735 35 9755 55
rect 9755 35 9760 55
rect 9730 30 9760 35
<< metal1 >>
rect 1670 13220 2000 13270
rect 1940 11340 2000 13220
rect 2540 11340 2580 11350
rect 1940 11300 2550 11340
rect 2570 11300 2580 11340
rect 2540 11290 2580 11300
rect 2140 11130 2180 11140
rect 2140 11110 2150 11130
rect 2170 11110 2180 11130
rect 2140 10750 2180 11110
rect 3580 11130 3620 11140
rect 3580 11110 3590 11130
rect 3610 11110 3620 11130
rect 3580 10750 3620 11110
rect 2140 10690 3620 10750
rect 2360 7940 2430 10690
rect 2770 10660 2820 10670
rect 2770 10640 2780 10660
rect 2810 10640 2820 10660
rect 2770 10630 2820 10640
rect 2770 10510 2810 10630
rect 2770 10480 2780 10510
rect 2800 10480 2810 10510
rect 2770 10470 2810 10480
rect 2040 7850 4380 7940
rect 4760 7850 6745 7940
rect 6855 7905 6965 7910
rect 6855 7885 6870 7905
rect 6940 7885 6965 7905
rect 6855 7875 6965 7885
rect 2040 7290 2080 7850
rect 2770 7750 2810 7780
rect 2770 7710 2780 7750
rect 2800 7710 2810 7750
rect 2770 7690 2810 7710
rect 2380 7340 2460 7350
rect 2380 7310 2390 7340
rect 2450 7310 2460 7340
rect 2380 7300 2460 7310
rect 2040 7270 2360 7290
rect 2040 7230 2300 7270
rect 2340 7230 2360 7270
rect 2040 7210 2360 7230
rect 1755 5210 1805 5220
rect 1755 5140 1765 5210
rect 1795 5180 1805 5210
rect 1795 5140 1810 5180
rect 1755 5130 1810 5140
rect 1620 5060 1805 5070
rect 1620 4990 1765 5060
rect 1795 5030 1805 5060
rect 1795 4990 1810 5030
rect 1620 4980 1810 4990
rect 1300 1460 1350 1480
rect 1300 1430 1310 1460
rect 1340 1430 1350 1460
rect 1300 820 1350 1430
rect -150 750 1350 820
rect 2040 830 2080 7210
rect 2380 7190 2460 7200
rect 2380 7160 2390 7190
rect 2450 7160 2460 7190
rect 2380 7070 2460 7160
rect 2380 6980 2480 7070
rect 2410 5330 2480 6980
rect 2770 5520 2805 7690
rect 2970 7595 6395 7695
rect 6300 6680 6395 7595
rect 6705 7275 6745 7850
rect 6705 6950 6750 7275
rect 6710 6865 6750 6950
rect 6930 6910 6965 7875
rect 7320 7005 7390 7015
rect 7320 6965 7340 7005
rect 7325 6935 7340 6965
rect 7370 6970 7390 7005
rect 7370 6940 7600 6970
rect 7370 6935 7385 6940
rect 7325 6930 7385 6935
rect 6930 6885 7465 6910
rect 6705 6855 7400 6865
rect 6705 6815 7200 6855
rect 6710 6810 6750 6815
rect 7185 6785 7200 6815
rect 7230 6815 7400 6855
rect 7230 6785 7245 6815
rect 7510 6800 7540 6875
rect 7185 6780 7245 6785
rect 7500 6785 7540 6800
rect 7500 6715 7505 6785
rect 7535 6715 7540 6785
rect 7500 6705 7540 6715
rect 6300 6590 7890 6680
rect 7555 5925 7635 6590
rect 7555 5825 7575 5925
rect 7615 5825 7635 5925
rect 7555 5810 7635 5825
rect 6980 5675 7745 5715
rect 8390 5675 8415 5680
rect 2765 5510 2815 5520
rect 2765 5440 2775 5510
rect 2805 5440 2815 5510
rect 2765 5430 2815 5440
rect 2410 5325 2735 5330
rect 6980 5325 7035 5675
rect 2410 5315 2950 5325
rect 2410 5295 2870 5315
rect 2940 5295 2950 5315
rect 2410 5285 2950 5295
rect 6800 5315 7035 5325
rect 6800 5295 6810 5315
rect 6880 5295 7035 5315
rect 6800 5285 7035 5295
rect 2410 2785 2485 5285
rect 2655 5210 2705 5220
rect 2655 5140 2665 5210
rect 2695 5180 2705 5210
rect 7320 5205 7390 5215
rect 7320 5180 7340 5205
rect 2695 5140 7340 5180
rect 2655 5135 7340 5140
rect 7370 5135 7390 5205
rect 2655 5130 7390 5135
rect 2655 5060 7610 5070
rect 2655 4990 2665 5060
rect 2695 5020 7610 5060
rect 2695 4990 2705 5020
rect 2655 4980 2705 4990
rect 7365 3620 7525 3645
rect 7365 3550 7480 3620
rect 7510 3550 7525 3620
rect 7365 3530 7525 3550
rect 7365 3350 7410 3530
rect 7570 3380 7610 5020
rect 8390 4955 8420 5675
rect 8400 3435 8430 3445
rect 8400 3410 8405 3435
rect 8425 3410 8430 3435
rect 8400 3400 8430 3410
rect 8500 3435 8680 3450
rect 8500 3410 8505 3435
rect 8525 3410 8680 3435
rect 8500 3400 8680 3410
rect 7185 3340 7245 3350
rect 7185 3270 7200 3340
rect 7230 3300 7245 3340
rect 7365 3325 7455 3350
rect 8400 3335 8430 3350
rect 8400 3310 8405 3335
rect 8425 3310 8430 3335
rect 8400 3300 8430 3310
rect 8500 3335 8560 3350
rect 8500 3310 8505 3335
rect 8525 3310 8560 3335
rect 8500 3300 8560 3310
rect 7230 3270 7455 3300
rect 7185 3255 7455 3270
rect 2410 2715 2430 2785
rect 2460 2715 2485 2785
rect 2410 2705 2485 2715
rect 2040 760 2050 830
rect 2070 760 2080 830
rect 2040 750 2080 760
rect 2190 2185 2875 2285
rect 2190 830 2255 2185
rect 2190 760 2205 830
rect 2225 760 2255 830
rect -150 550 -70 750
rect 2190 745 2255 760
rect 2415 2125 2800 2150
rect 2415 2055 2430 2125
rect 2460 2055 2800 2125
rect 2415 2050 2800 2055
rect 7500 2120 7790 2150
rect 2415 655 2480 2050
rect 7500 1000 7560 2120
rect 7500 970 7510 1000
rect 7540 970 7560 1000
rect 7500 960 7560 970
rect 0 570 10 640
rect 2040 560 2480 655
rect -3100 540 -70 550
rect -3100 520 -3090 540
rect -3070 520 -2670 540
rect -2650 520 -2220 540
rect -2200 520 -1770 540
rect -1750 520 -1320 540
rect -1300 520 -900 540
rect -880 520 -450 540
rect -430 520 -70 540
rect -3100 510 -70 520
rect -3100 270 -100 280
rect -3100 250 -3090 270
rect -3070 250 -2670 270
rect -2650 250 -2220 270
rect -2200 250 -1770 270
rect -1750 250 -1320 270
rect -1300 250 -900 270
rect -880 250 -450 270
rect -430 250 -100 270
rect -3100 240 -100 250
rect -150 50 -100 240
rect 2755 80 2820 90
rect -150 0 620 50
rect 570 -30 620 0
rect 940 0 1010 40
rect 2755 20 2775 80
rect 2040 10 2775 20
rect 2805 60 2820 80
rect 2805 45 2920 60
rect 2805 25 2840 45
rect 2910 25 2920 45
rect 2805 10 2920 25
rect 2040 0 2920 10
rect 8520 10 8560 3300
rect 8640 1380 8680 3400
rect 8640 1320 9840 1380
rect 9180 1260 9230 1270
rect 9180 1230 9190 1260
rect 9220 1230 9230 1260
rect 9180 60 9230 1230
rect 9790 410 9840 1320
rect 9790 380 9800 410
rect 9830 380 9840 410
rect 9790 370 9840 380
rect 9180 30 9190 60
rect 9220 30 9230 60
rect 9180 20 9230 30
rect 9720 60 9770 70
rect 9720 30 9730 60
rect 9760 30 9770 60
rect 9720 10 9770 30
rect 8520 0 9160 10
rect 9260 0 9770 10
rect 940 -30 980 0
rect 8520 -30 9770 0
rect 570 -70 980 -30
<< via1 >>
rect 1765 5140 1795 5210
rect 1765 4990 1795 5060
rect 7340 6935 7370 7005
rect 7200 6785 7230 6855
rect 7505 6715 7535 6785
rect 7575 5825 7615 5925
rect 2775 5440 2805 5510
rect 2665 5140 2695 5210
rect 7340 5135 7370 5205
rect 2665 4990 2695 5060
rect 7480 3550 7510 3620
rect 7200 3270 7230 3340
rect 7945 3040 7975 3110
rect 2430 2715 2460 2785
rect 2430 2055 2460 2125
rect 2775 10 2805 80
<< metal2 >>
rect 7325 7005 7385 7015
rect 7325 6970 7340 7005
rect 7320 6935 7340 6970
rect 7370 6935 7385 7005
rect 7320 6930 7385 6935
rect 7185 6855 7245 6865
rect 7185 6785 7200 6855
rect 7230 6785 7245 6855
rect 2765 5510 2815 5520
rect 2765 5440 2775 5510
rect 2805 5440 2815 5510
rect 1650 5210 2710 5220
rect 1650 5140 1765 5210
rect 1795 5140 2665 5210
rect 2695 5140 2710 5210
rect 1650 5130 2710 5140
rect 1750 5060 2710 5070
rect 1750 4990 1765 5060
rect 1795 4990 2665 5060
rect 2695 4990 2710 5060
rect 1750 4980 2710 4990
rect 2420 2785 2470 2805
rect 2420 2715 2430 2785
rect 2460 2715 2470 2785
rect 2420 2125 2470 2715
rect 2420 2055 2430 2125
rect 2460 2055 2470 2125
rect 2420 2045 2470 2055
rect 2765 80 2815 5440
rect 7185 3340 7245 6785
rect 7320 5215 7380 6930
rect 7500 6785 7540 6800
rect 7500 6715 7505 6785
rect 7535 6715 7540 6785
rect 7320 5210 7385 5215
rect 7325 5205 7385 5210
rect 7325 5135 7340 5205
rect 7370 5135 7385 5205
rect 7325 5130 7385 5135
rect 7500 3640 7540 6715
rect 7555 5925 7635 5970
rect 7555 5825 7575 5925
rect 7615 5825 7635 5925
rect 7555 5810 7635 5825
rect 7560 4460 7635 5810
rect 7560 4390 7645 4460
rect 7560 4385 7940 4390
rect 7560 4280 7995 4385
rect 7465 3620 7540 3640
rect 7465 3550 7480 3620
rect 7510 3550 7540 3620
rect 7465 3535 7540 3550
rect 7185 3270 7200 3340
rect 7230 3270 7245 3340
rect 7185 3260 7245 3270
rect 7920 3110 7995 4280
rect 7920 3040 7945 3110
rect 7975 3040 7995 3110
rect 7920 3010 7995 3040
rect 2765 10 2775 80
rect 2805 10 2815 80
rect 2765 0 2815 10
use bbg  bbg_0
timestamp 1762117721
transform 1 0 220 0 1 560
box -220 -560 1820 210
use ccm  ccm_0
timestamp 1762197520
transform 1 0 9265 0 1 25
box -1810 -10 2910 1120
use dac  dac_0
timestamp 1762200396
transform 1 0 -2430 0 1 9720
box -620 -8740 4340 3870
use fvf  fvf_0
timestamp 1762117721
transform 0 1 7910 -1 0 8390
box -150 -510 3125 510
use fvf  fvf_1
timestamp 1762117721
transform 0 1 7960 -1 0 4830
box -150 -510 3125 510
use inv  inv_0
timestamp 1762200811
transform 1 0 -380 0 1 160
box -90 -50 200 490
use inv  inv_1
timestamp 1762200811
transform 1 0 -830 0 1 160
box -90 -50 200 490
use inv  inv_2
timestamp 1762200811
transform 1 0 -1250 0 1 160
box -90 -50 200 490
use inv  inv_3
timestamp 1762200811
transform 1 0 -1700 0 1 160
box -90 -50 200 490
use inv  inv_4
timestamp 1762200811
transform 1 0 -3020 0 1 160
box -90 -50 200 490
use inv  inv_6
timestamp 1762200811
transform 1 0 -2600 0 1 160
box -90 -50 200 490
use inv  inv_7
timestamp 1762200811
transform 1 0 -2150 0 1 160
box -90 -50 200 490
use ncbc  ncbc_0
timestamp 1762137910
transform 1 0 3155 0 1 4445
box -350 810 3735 5830
use pcbc  pcbc_0
timestamp 1762135317
transform 1 0 -1317 0 1 -2702
box 4115 2710 8150 7690
<< labels >>
rlabel locali 9745 25 9745 25 5 Vcn
port 3 s
<< end >>
