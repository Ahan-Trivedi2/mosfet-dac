* SPICE3 file created from full.ext - technology: sky130A

.subckt dac Iout Idump VN Iin Vg b6 bn6 b5 bn5 b4 bn4 b3 bn3 b2 bn2 b1 bn1 b0 bn0
X0 a_6220_2110# b0 a_6220_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X1 a_2270_n1450# Vg a_2270_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X2 a_3350_n7120# Vg a_3350_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X3 a_1900_3210# b4 a_1900_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X4 a_4060_n7120# Vg a_4060_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X5 VN VN Idump VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X6 a_110_n350# Vg a_110_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X7 VN VN a_3350_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X8 a_3350_n2550# Vg a_2270_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X9 VN VN a_4430_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X10 a_4060_n2550# Vg a_3350_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X11 a_4430_n8220# Vg a_4430_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X12 a_5140_n8220# Vg a_5140_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X13 a_5140_4310# b1 a_5140_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X14 a_4060_n10730# b2 a_4060_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X15 a_4430_3210# bn2 a_4430_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X16 a_3350_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X17 a_n260_n9320# Vg a_n260_n10730# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X18 a_4430_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X19 VN VN a_110_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X20 a_1190_n10420# Vg a_1900_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X21 a_4060_n14030# b2 Iout VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X22 a_5140_n11830# b1 a_5140_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X23 a_6220_n10730# bn0 a_6590_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X24 VN VN Idump VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X25 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X26 a_820_n8220# Vg a_820_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X27 Iout VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X28 a_2270_n9320# Vg a_2270_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X29 a_4430_n350# Vg a_4430_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X30 a_1900_n1450# Vg a_1900_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X31 a_6590_n14030# bn0 Idump VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X32 a_6220_n12930# b0 a_6220_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X33 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X34 a_5140_n350# Vg a_5140_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X35 a_2270_n10420# Vg a_2980_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X36 a_4430_n10420# Vg a_5510_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X37 a_1900_n12930# b4 a_1900_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X38 Idump bn3 a_3350_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X39 a_3350_750# Vg a_3350_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X40 a_110_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X41 a_5510_n10420# Vg a_6220_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X42 a_110_3210# bn6 a_110_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X43 a_820_3210# b5 a_820_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X44 a_2980_n1450# Vg a_2980_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X45 a_5510_n1450# Vg a_5510_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X46 a_4060_3210# b2 a_4060_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X47 a_6220_n1450# Vg a_6220_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X48 a_5510_n10420# Vg a_6590_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X49 a_7300_n7120# Vg a_7300_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X50 a_3350_2110# bn3 a_2980_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X51 a_820_n350# Vg a_820_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X52 a_n260_n11830# b6 a_n260_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X53 Idump bn0 a_6590_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X54 a_6590_750# Vg a_6590_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X55 a_820_n10730# bn5 a_1190_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X56 a_6590_n1450# Vg a_6590_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X57 a_7300_n2550# Vg a_6590_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X58 Iout VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X59 a_1190_n14030# bn5 Idump VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X60 a_2270_n11830# bn4 a_2270_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X61 a_6590_2110# bn0 a_6220_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X62 VN VN Iin VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X63 a_5510_n9320# Vg a_5510_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X64 a_2270_4310# bn4 a_2270_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X65 a_2980_4310# b3 a_2980_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X66 Idump VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X67 a_3350_n12930# bn3 a_3350_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X68 a_n260_n8220# Vg a_n260_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X69 a_110_n12930# bn6 a_110_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X70 Iin VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X71 VN VN Idump VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X72 a_4060_n10730# bn2 a_4430_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X73 a_820_n9320# Vg a_820_n10730# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X74 Idump Vg a_7300_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X75 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X76 a_n260_n350# Vg a_n260_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X77 a_4430_n14030# bn2 Idump VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X78 a_5510_n11830# bn1 a_5510_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X79 a_1190_3210# bn5 a_1190_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X80 a_1190_n7120# Vg a_1190_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X81 a_2980_n10730# b3 a_2980_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X82 VN VN a_1190_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X83 Idump VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X84 a_n260_3210# b6 a_n260_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X85 a_2980_n14030# b3 Iout VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X86 VN VN Idump VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X87 a_1190_n2550# Vg a_110_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X88 a_2270_n8220# Vg a_2270_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X89 a_110_n7120# Vg a_110_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X90 a_820_n11830# b5 a_820_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X91 a_6220_4310# b0 a_6220_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X92 a_5510_3210# bn1 a_5510_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X93 a_1190_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X94 Iout b4 a_1900_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X95 a_1900_750# Vg a_1900_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X96 a_110_n2550# Vg Iin VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X97 Iout VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X98 a_2270_n350# Vg a_2270_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X99 a_2270_n10420# Vg a_3350_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X100 a_1900_2110# b4 a_1900_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X101 a_3350_n10420# Vg a_4060_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X102 a_6220_n9320# Vg a_6220_n10730# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X103 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X104 Idump bn2 a_4430_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X105 VN VN a_1190_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X106 a_4060_n12930# b2 a_4060_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X107 a_1900_n9320# Vg a_1900_n10730# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X108 a_4430_750# Vg a_4430_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X109 a_3350_n1450# Vg a_3350_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X110 a_4060_n1450# Vg a_4060_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X111 a_4430_n7120# Vg a_4430_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X112 a_1900_n8220# Vg a_1900_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X113 a_5140_n7120# Vg a_5140_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X114 a_6590_n12930# bn0 a_6590_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X115 a_5140_3210# b1 a_5140_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X116 VN VN a_2270_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X117 VN VN a_4430_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X118 VN VN a_5510_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X119 a_4430_2110# bn2 a_4060_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X120 a_4430_n2550# Vg a_3350_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X121 a_1190_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X122 a_5140_n2550# Vg a_4430_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X123 a_5140_n10730# b1 a_5140_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X124 a_5510_n8220# Vg a_5510_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X125 a_2980_n8220# Vg a_2980_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X126 a_6220_n8220# Vg a_6220_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X127 Idump bn6 a_110_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X128 Iout b5 a_820_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X129 a_110_750# Vg a_110_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X130 a_820_750# Vg a_820_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X131 VN VN a_5510_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X132 a_820_n7120# Vg a_820_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X133 a_1900_n350# Vg a_1900_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X134 a_2270_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X135 a_4430_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X136 a_5140_n14030# b1 Iout VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X137 a_6220_n11830# b0 a_6220_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X138 Iout b2 a_4060_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X139 a_4060_750# Vg a_4060_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X140 a_5510_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X141 a_1900_n11830# b4 a_1900_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X142 a_6590_n8220# Vg a_6590_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X143 a_3350_4310# bn3 a_3350_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X144 a_820_n2550# Vg a_110_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X145 Iout VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X146 a_3350_n9320# Vg a_3350_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X147 a_110_2110# bn6 a_n260_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X148 a_820_2110# b5 a_820_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X149 Iout VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X150 a_1190_n12930# bn5 a_1190_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X151 a_2980_n350# Vg a_2980_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X152 a_5510_n350# Vg a_5510_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X153 a_5510_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X154 a_4060_2110# b2 a_4060_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X155 a_6220_n350# Vg a_6220_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X156 a_110_n9320# Vg a_110_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X157 a_6590_n10420# Vg a_7300_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X158 a_n260_n10730# b6 a_n260_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X159 a_6590_4310# bn0 a_6590_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X160 VN VN Idump VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X161 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X162 a_6590_n350# Vg a_6590_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X163 a_7300_n1450# Vg a_7300_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X164 a_n260_n14030# b6 Iout VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X165 a_1900_n10730# bn4 a_2270_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X166 a_2270_3210# bn4 a_2270_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X167 a_2980_3210# b3 a_2980_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X168 a_2270_n14030# bn4 Idump VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X169 a_3350_n11830# bn3 a_3350_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X170 a_n260_n7120# Vg a_n260_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X171 Idump VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X172 a_4430_n12930# bn2 a_4430_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X173 a_110_n11830# bn6 a_110_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X174 a_n260_n2550# Vg Iin VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X175 Idump bn5 a_1190_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X176 a_1190_750# Vg a_1190_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X177 Idump VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X178 a_2980_n12930# b3 a_2980_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X179 Iout b6 a_n260_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X180 a_n260_750# Vg a_n260_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X181 a_5140_n10730# bn1 a_5510_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X182 a_1190_2110# bn5 a_820_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X183 a_110_n10420# Vg a_1190_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X184 a_5510_n14030# bn1 Idump VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X185 a_n260_2110# b6 a_n260_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X186 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X187 Idump bn1 a_5510_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X188 a_1190_n1450# Vg a_1190_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X189 a_4060_n9320# Vg a_4060_n10730# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X190 a_5510_750# Vg a_5510_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X191 a_2270_n7120# Vg a_2270_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X192 VN VN a_2270_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X193 a_6590_n9320# Vg a_6590_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X194 VN VN a_3350_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X195 Iin Vg a_110_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X196 a_820_n10730# b5 a_820_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X197 a_6220_3210# b0 a_6220_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X198 a_5510_2110# bn1 a_5140_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X199 a_2270_n2550# Vg a_1190_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X200 a_3350_n8220# Vg a_3350_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X201 a_1900_4310# b4 a_1900_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X202 a_820_n14030# b5 Iout VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X203 a_4060_n8220# Vg a_4060_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X204 a_110_n1450# Vg a_110_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X205 a_2270_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X206 a_3350_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X207 Iout b1 a_5140_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X208 a_5140_750# Vg a_5140_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X209 a_4060_n11830# b2 a_4060_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X210 a_4430_4310# bn2 a_4430_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X211 a_7300_n9320# Vg Idump VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X212 a_3350_n350# Vg a_3350_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X213 a_4060_n350# Vg a_4060_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X214 a_3350_n10420# Vg a_4430_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X215 a_1900_n7120# Vg a_1900_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X216 Iout VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X217 a_5140_n12930# b1 a_5140_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X218 a_1190_n9320# Vg a_1190_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X219 a_4430_n10420# Vg a_5140_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X220 a_6590_n11830# bn0 a_6590_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X221 a_5140_2110# b1 a_5140_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X222 a_4430_n1450# Vg a_4430_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X223 a_1900_n2550# Vg a_1190_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X224 Idump VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X225 a_5140_n1450# Vg a_5140_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X226 a_2980_n7120# Vg a_2980_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X227 a_5510_n7120# Vg a_5510_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X228 VN VN Idump VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X229 a_6220_n7120# Vg a_6220_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X230 a_110_4310# bn6 a_110_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X231 a_820_4310# b5 a_820_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X232 VN VN a_6590_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X233 a_110_n10420# Vg a_820_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X234 a_2980_n2550# Vg a_2270_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X235 a_5510_n2550# Vg a_4430_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X236 a_6220_n10730# b0 a_6220_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X237 a_4060_4310# b2 a_4060_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X238 a_6220_n2550# Vg a_5510_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X239 a_6590_n7120# Vg a_6590_n8220# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X240 a_1900_n10730# b4 a_1900_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X241 a_7300_n8220# Vg a_7300_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X242 a_3350_3210# bn3 a_3350_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X243 a_820_n1450# Vg a_820_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X244 a_6220_n14030# b0 Iout VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X245 a_n260_n12930# b6 a_n260_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X246 VN VN Idump VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X247 a_1900_n14030# b4 Iout VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X248 a_1190_n11830# bn5 a_1190_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X249 a_6590_n2550# Vg a_5510_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X250 a_6590_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X251 a_4430_n9320# Vg a_4430_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X252 Idump VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X253 a_2270_n12930# bn4 a_2270_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X254 a_6590_3210# bn0 a_6590_2110# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X255 a_2980_n9320# Vg a_2980_n10730# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X256 Idump bn4 a_2270_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X257 Iout b3 a_2980_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X258 a_2270_750# Vg a_2270_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X259 a_2980_750# Vg a_2980_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X260 a_7300_n350# Vg a_7300_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X261 a_2270_2110# bn4 a_1900_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X262 a_2980_2110# b3 a_2980_750# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X263 a_2980_n10730# bn3 a_3350_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X264 Iin Vg a_n260_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X265 a_3350_n14030# bn3 Idump VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X266 a_4430_n11830# bn2 a_4430_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X267 VN VN a_110_n10420# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X268 Idump VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X269 a_n260_n10730# bn6 a_110_n11830# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X270 a_n260_n1450# Vg a_n260_n2550# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X271 a_5510_n12930# bn1 a_5510_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X272 a_1190_4310# bn5 a_1190_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X273 a_1190_n8220# Vg a_1190_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X274 a_110_n14030# bn6 Idump VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X275 a_2980_n11830# b3 a_2980_n12930# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X276 a_n260_4310# b6 a_n260_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X277 Iout VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X278 a_110_750# VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X279 VN VN Iin VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X280 a_110_n8220# Vg a_110_n9320# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X281 a_820_n12930# b5 a_820_n14030# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X282 Iout b0 a_6220_4310# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X283 a_5510_4310# bn1 a_5510_3210# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X284 a_6220_750# Vg a_6220_n350# VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X285 a_1190_n350# Vg a_1190_n1450# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X286 VN VN Iout VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X287 Iin VN VN VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X288 a_1190_n10420# Vg a_2270_n7120# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X289 a_5140_n9320# Vg a_5140_n10730# VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
.ends

.subckt pcbc VN Vbn Vc VP
X0 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X1 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X2 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X3 a_8360_6840# a_8320_6920# VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X4 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X5 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X6 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X7 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X8 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X9 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X10 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X11 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X12 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X13 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X14 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X15 a_8360_6840# a_8320_6920# VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X16 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X17 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X18 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X19 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X20 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X21 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X22 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X23 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X24 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X25 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X26 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X27 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X28 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X29 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X30 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X31 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X32 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X33 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X34 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X35 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X36 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X37 VP a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X38 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X39 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X40 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X41 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X42 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X43 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X44 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X45 Vc Vc a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X46 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X47 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X48 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X49 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X50 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X51 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X52 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X53 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X54 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X55 Vc Vc a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X56 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X57 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X58 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X59 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X60 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X61 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X62 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X63 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X64 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X65 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X66 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X67 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X68 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X69 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X70 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X71 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X72 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X73 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X74 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X75 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X76 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X77 a_8360_6840# Vc Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X78 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X79 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X80 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X81 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X82 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X83 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X84 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X85 VP VP a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X86 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X87 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X88 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X89 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X90 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X91 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X92 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X93 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X94 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X95 VP VP a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X96 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X97 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X98 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X99 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X100 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X101 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X102 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X103 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X104 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X105 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X106 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X107 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X108 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X109 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X110 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X111 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X112 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X113 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X114 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X115 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X116 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X117 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X118 a_8360_6840# VP VP VP sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X119 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X120 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X121 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X122 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X123 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X124 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X125 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X126 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X127 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X128 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X129 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X130 VP a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X131 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X132 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X133 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X134 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X135 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X136 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X137 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X138 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X139 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X140 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X141 a_8360_6840# VP VP VP sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X142 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X143 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X144 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X145 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X146 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X147 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X148 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X149 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X150 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X151 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X152 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X153 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X154 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X155 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X156 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X157 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X158 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X159 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X160 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X161 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X162 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X163 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X164 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X165 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X166 a_8360_6840# Vc Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X167 a_8320_6920# a_8320_6920# a_8360_6840# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X168 a_8360_6840# a_8320_6920# a_8320_6920# VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X169 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X170 VN Vbn a_8320_6920# VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X171 a_8320_6920# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
.ends

.subckt ccm VP VN Vdsg Vcn Vcp Vout
X0 VP a_3280_100# a_3480_1180# VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X1 a_3280_100# Vcn a_2200_100# VN sky130_fd_pr__nfet_01v8 ad=0.87 pd=5.3 as=0.58 ps=3.53 w=2 l=5
X2 a_2200_100# Vdsg VN VN sky130_fd_pr__nfet_01v8 ad=0.58 pd=3.53 as=2.14 ps=7 w=2 l=5
X3 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=24.6 ps=113.2 w=2 l=5
X4 Vout VP VP VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=1.47 ps=5.9 w=2 l=5
X5 VP a_3280_100# a_3280_100# VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.87 ps=5.3 w=2 l=5
X6 Vout VP VP VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=1.47 ps=5.9 w=2 l=5
X7 VN Vdsg a_n80_100# VN sky130_fd_pr__nfet_01v8 ad=2.14 pd=7 as=0.58 ps=3.53 w=2 l=5
X8 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0 ps=0 w=2 l=5
X9 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0 ps=0 w=2 l=5
X10 Vout Vcp a_n1360_1180# VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X11 Vout Vcp a_n1360_1180# VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X12 VP VP Vout VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0.58 ps=3.53 w=2 l=5
X13 VP VP Vout VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0.58 ps=3.53 w=2 l=5
X14 a_2200_100# Vdsg VN VN sky130_fd_pr__nfet_01v8 ad=0.58 pd=3.53 as=2.14 ps=7 w=2 l=5
X15 a_n80_100# Vcn a_n2360_60# VN sky130_fd_pr__nfet_01v8 ad=0.58 pd=3.53 as=0.87 ps=5.3 w=2 l=5
X16 VN Vdsg a_n80_100# VN sky130_fd_pr__nfet_01v8 ad=2.14 pd=7 as=0.58 ps=3.53 w=2 l=5
X17 a_n1360_1180# a_n2360_60# VP VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X18 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0 ps=0 w=2 l=5
X19 a_n1360_1180# a_n2360_60# VP VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X20 a_n2360_60# a_n2360_60# VP VP sky130_fd_pr__pfet_01v8 ad=0.87 pd=5.3 as=0.58 ps=3.53 w=2 l=5
X21 a_n80_100# Vcn a_n2360_60# VN sky130_fd_pr__nfet_01v8 ad=0.58 pd=3.53 as=0.87 ps=5.3 w=2 l=5
X22 a_3480_1180# Vcp Vout VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X23 a_3480_1180# Vcp Vout VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X24 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0 ps=0 w=2 l=5
X25 a_3280_100# Vcn a_2200_100# VN sky130_fd_pr__nfet_01v8 ad=0.87 pd=5.3 as=0.58 ps=3.53 w=2 l=5
X26 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0 ps=0 w=2 l=5
X27 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0 ps=0 w=2 l=5
X28 a_n2360_60# a_n2360_60# VP VP sky130_fd_pr__pfet_01v8 ad=0.87 pd=5.3 as=0.58 ps=3.53 w=2 l=5
X29 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0 ps=0 w=2 l=5
X30 VP a_3280_100# a_3480_1180# VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X31 VP a_3280_100# a_3280_100# VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.87 ps=5.3 w=2 l=5
.ends

.subckt inv A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.5
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.5
X2 VP A Y VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5
X3 VN A Y VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5
.ends

.subckt ncbc Vc Vp Vbp Vn
X0 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X1 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X2 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X3 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X4 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X5 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X6 a_n560_3080# Vc Vc Vn sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X7 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X8 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X9 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X10 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X11 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X12 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X13 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X14 Vc Vc a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X15 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X16 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X17 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X18 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X19 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X20 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X21 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X22 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X23 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X24 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X25 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X26 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X27 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X28 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X29 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X30 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X31 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X32 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X33 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X34 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X35 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X36 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X37 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X38 Vc Vc a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X39 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X40 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X41 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X42 a_n560_3080# Vn Vn Vn sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X43 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X44 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X45 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X46 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X47 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X48 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X49 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X50 Vn a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X51 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X52 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X53 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X54 a_n560_3080# a_n600_3160# Vn Vn sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X55 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X56 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X57 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X58 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X59 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X60 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X61 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X62 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X63 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X64 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X65 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X66 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X67 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X68 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X69 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X70 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X71 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X72 Vn Vn a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X73 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X74 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X75 a_n560_3080# Vc Vc Vn sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X76 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X77 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X78 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X79 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X80 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X81 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X82 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X83 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X84 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X85 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X86 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X87 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X88 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X89 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X90 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X91 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X92 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X93 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X94 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X95 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X96 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X97 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X98 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X99 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X100 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X101 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X102 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X103 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X104 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X105 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X106 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X107 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X108 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X109 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X110 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X111 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X112 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X113 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X114 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X115 Vn a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X116 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X117 a_n560_3080# a_n600_3160# Vn Vn sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X118 a_n560_3080# Vn Vn Vn sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X119 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X120 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X121 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X122 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X123 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X124 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X125 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X126 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X127 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X128 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X129 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X130 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X131 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X132 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X133 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X134 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X135 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X136 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X137 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X138 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X139 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X140 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X141 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X142 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X143 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X144 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X145 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X146 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X147 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X148 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X149 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X150 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X151 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X152 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X153 Vn Vn a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X154 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X155 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X156 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X157 a_n600_3160# a_n600_3160# a_n560_3080# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X158 Vp Vp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X159 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X160 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X161 Vp Vbp a_n600_3160# Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X162 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X163 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X164 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X165 a_n600_3160# Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X166 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X167 Vp Vbp Vc Vp sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X168 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X169 a_n560_3080# a_n600_3160# a_n600_3160# Vn sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X170 Vc Vp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X171 Vc Vbp Vp Vp sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
.ends

.subckt bbg VP VBP VBN VN RES
X0 VN a_460_n780# a_n200_n840# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X1 a_460_n780# VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X2 a_460_n780# a_460_n780# RES VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X3 VP VBP a_460_n780# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X4 a_n200_n840# a_460_n780# VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X5 VP a_n200_n840# a_n200_n840# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X6 VN VBN VBP VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X7 VBP a_n200_n840# VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X8 VBN VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X9 a_n200_n840# a_460_n780# VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X10 RES a_460_n780# a_460_n780# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X11 VP VBP VBN VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X12 VP VBP VBN VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X13 VBP a_n200_n840# VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X14 a_n200_n840# a_n200_n840# VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X15 VBP VBN VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X16 a_460_n780# VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X17 a_460_n780# a_460_n780# RES VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X18 VP VBP a_460_n780# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X19 VBN VBN VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X20 VBN VBN VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X21 VP a_n200_n840# a_n200_n840# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X22 VN VBN VBP VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X23 RES a_460_n780# a_460_n780# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X24 VN VBN VBN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X25 VP a_n200_n840# VBP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X26 VP a_n200_n840# VBP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X27 VN VBN VBN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X28 VN a_460_n780# a_n200_n840# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X29 VBP VBN VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X30 VBN VBP VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X31 a_n200_n840# a_n200_n840# VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
.ends

.subckt fvf VP Vdsg VN Vin Vc Vbp
X0 Vin Vc Vdsg VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=1 ps=5 w=2 l=5
X1 Vin Vdsg VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=5
X2 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=4 ps=24 w=1 l=1
X3 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=1
X4 Vdsg Vc Vin VN sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0.5 ps=2.5 w=2 l=5
X5 Vdsg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=1
X6 Vin Vc Vdsg VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=1 ps=5 w=2 l=5
X7 VP Vbp Vdsg VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1
X8 Vdsg Vc Vin VN sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0.5 ps=2.5 w=2 l=5
X9 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=1
X10 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=1
X11 VN Vdsg Vin VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=5
X12 Vin Vdsg VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=5
X13 Vdsg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=1
X14 VP Vbp Vdsg VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1
X15 VN Vdsg Vin VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=5
.ends

.subckt full Vcn
Xdac_0 fvf_1/Vin fvf_0/Vin Vcn dac_0/Iin inv_7/VP inv_4/A inv_4/Y inv_6/A inv_6/Y
+ inv_7/A inv_7/Y inv_3/A inv_3/Y inv_2/A inv_2/Y inv_1/A inv_1/Y inv_0/A inv_0/Y
+ dac
Xpcbc_0 Vcn bbg_0/VBN pcbc_0/Vc fvf_1/VP pcbc
Xccm_0 fvf_1/VP Vcn Vcn fvf_1/Vc pcbc_0/Vc ccm_0/Vout ccm
Xinv_0 inv_0/A inv_0/Y inv_7/VP Vcn inv
Xinv_1 inv_1/A inv_1/Y inv_7/VP Vcn inv
Xinv_2 inv_2/A inv_2/Y inv_7/VP Vcn inv
Xinv_3 inv_3/A inv_3/Y inv_7/VP Vcn inv
Xinv_4 inv_4/A inv_4/Y inv_7/VP Vcn inv
Xncbc_0 fvf_1/Vc fvf_1/VP fvf_1/Vbp Vcn ncbc
Xinv_7 inv_7/A inv_7/Y inv_7/VP Vcn inv
Xinv_6 inv_6/A inv_6/Y inv_7/VP Vcn inv
Xbbg_0 fvf_1/VP fvf_1/Vbp bbg_0/VBN Vcn bbg_0/RES bbg
Xfvf_0 fvf_1/VP fvf_0/Vdsg Vcn fvf_0/Vin fvf_1/Vc fvf_1/Vbp fvf
Xfvf_1 fvf_1/VP Vcn Vcn fvf_1/Vin fvf_1/Vc fvf_1/Vbp fvf
X0 Vcn a_5360_22280# a_5360_22280# Vcn sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=1
X1 inv_7/VP fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=3
X2 a_5360_22280# a_5360_22280# Vcn Vcn sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=1
X3 fvf_1/VP fvf_1/Vbp inv_7/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=3
X4 a_5360_22280# inv_7/VP inv_7/VP Vcn sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=1
X5 inv_7/VP inv_7/VP a_5360_22280# Vcn sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=1
X6 a_5360_22280# a_5360_22280# Vcn Vcn sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=1
X7 Vcn a_5360_22280# a_5360_22280# Vcn sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=1
X8 inv_7/VP inv_7/VP a_5360_22280# Vcn sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=1
X9 a_5360_22280# inv_7/VP inv_7/VP Vcn sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=1
X10 inv_7/VP fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=3
X11 fvf_1/VP fvf_1/Vbp inv_7/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=3
X12 dac_0/Iin fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
.ends

