magic
tech sky130A
timestamp 1762049146
<< nwell >>
rect -330 5270 -90 6630
rect 3410 5270 3650 6630
rect -330 4910 3650 5270
rect -330 3550 -90 4910
rect 3410 3550 3650 4910
<< nmos >>
rect -30 6610 70 7610
rect 140 6610 240 7610
rect 310 6610 410 7610
rect 480 6610 580 7610
rect 650 6610 750 7610
rect 820 6610 920 7610
rect 990 6610 1090 7610
rect 1160 6610 1260 7610
rect 1330 6610 1430 7610
rect 1500 6610 1600 7610
rect 1720 6610 1820 7610
rect 1890 6610 1990 7610
rect 2060 6610 2160 7610
rect 2230 6610 2330 7610
rect 2400 6610 2500 7610
rect 2570 6610 2670 7610
rect 2740 6610 2840 7610
rect 2910 6610 3010 7610
rect 3080 6610 3180 7610
rect 3250 6610 3350 7610
rect -30 5570 70 6570
rect 140 5570 240 6570
rect 310 5570 410 6570
rect 480 5570 580 6570
rect 650 5570 750 6570
rect 820 5570 920 6570
rect 990 5570 1090 6570
rect 1160 5570 1260 6570
rect 1330 5570 1430 6570
rect 1500 5570 1600 6570
rect -30 5360 70 5460
rect 140 5360 240 5460
rect 310 5360 410 5460
rect 480 5360 580 5460
rect 650 5360 750 5460
rect 820 5360 920 5460
rect 990 5360 1090 5460
rect 1160 5360 1260 5460
rect 1330 5360 1430 5460
rect 1500 5360 1600 5460
rect 1720 5570 1820 6570
rect 1890 5570 1990 6570
rect 2060 5570 2160 6570
rect 2230 5570 2330 6570
rect 2400 5570 2500 6570
rect 2570 5570 2670 6570
rect 2740 5570 2840 6570
rect 2910 5570 3010 6570
rect 3080 5570 3180 6570
rect 3250 5570 3350 6570
rect 1720 5360 1820 5460
rect 1890 5360 1990 5460
rect 2060 5360 2160 5460
rect 2230 5360 2330 5460
rect 2400 5360 2500 5460
rect 2570 5360 2670 5460
rect 2740 5360 2840 5460
rect 2910 5360 3010 5460
rect 3080 5360 3180 5460
rect 3250 5360 3350 5460
rect -30 4720 70 4820
rect 140 4720 240 4820
rect 310 4720 410 4820
rect 480 4720 580 4820
rect 650 4720 750 4820
rect 820 4720 920 4820
rect 990 4720 1090 4820
rect 1160 4720 1260 4820
rect 1330 4720 1430 4820
rect 1500 4720 1600 4820
rect -30 3610 70 4610
rect 140 3610 240 4610
rect 310 3610 410 4610
rect 480 3610 580 4610
rect 650 3610 750 4610
rect 820 3610 920 4610
rect 990 3610 1090 4610
rect 1160 3610 1260 4610
rect 1330 3610 1430 4610
rect 1500 3610 1600 4610
rect 1720 4720 1820 4820
rect 1890 4720 1990 4820
rect 2060 4720 2160 4820
rect 2230 4720 2330 4820
rect 2400 4720 2500 4820
rect 2570 4720 2670 4820
rect 2740 4720 2840 4820
rect 2910 4720 3010 4820
rect 3080 4720 3180 4820
rect 3250 4720 3350 4820
rect 1720 3610 1820 4610
rect 1890 3610 1990 4610
rect 2060 3610 2160 4610
rect 2230 3610 2330 4610
rect 2400 3610 2500 4610
rect 2570 3610 2670 4610
rect 2740 3610 2840 4610
rect 2910 3610 3010 4610
rect 3080 3610 3180 4610
rect 3250 3610 3350 4610
rect -30 2570 70 3570
rect 140 2570 240 3570
rect 310 2570 410 3570
rect 480 2570 580 3570
rect 650 2570 750 3570
rect 820 2570 920 3570
rect 990 2570 1090 3570
rect 1160 2570 1260 3570
rect 1330 2570 1430 3570
rect 1500 2570 1600 3570
rect 1720 2570 1820 3570
rect 1890 2570 1990 3570
rect 2060 2570 2160 3570
rect 2230 2570 2330 3570
rect 2400 2570 2500 3570
rect 2570 2570 2670 3570
rect 2740 2570 2840 3570
rect 2910 2570 3010 3570
rect 3080 2570 3180 3570
rect 3250 2570 3350 3570
<< pmos >>
rect -310 6070 -110 6570
rect -310 5530 -110 6030
rect 3430 6070 3630 6570
rect 3430 5530 3630 6030
rect -190 5140 -90 5240
rect -50 5140 50 5240
rect 90 5140 190 5240
rect 230 5140 330 5240
rect 370 5140 470 5240
rect 510 5140 610 5240
rect 650 5140 750 5240
rect 790 5140 890 5240
rect 930 5140 1030 5240
rect 1070 5140 1170 5240
rect 1210 5140 1310 5240
rect 2010 5140 2110 5240
rect 2150 5140 2250 5240
rect 2290 5140 2390 5240
rect 2430 5140 2530 5240
rect 2570 5140 2670 5240
rect 2710 5140 2810 5240
rect 2850 5140 2950 5240
rect 2990 5140 3090 5240
rect 3130 5140 3230 5240
rect 3270 5140 3370 5240
rect 3410 5140 3510 5240
rect -190 4940 -90 5040
rect -50 4940 50 5040
rect 90 4940 190 5040
rect 230 4940 330 5040
rect 370 4940 470 5040
rect 510 4940 610 5040
rect 650 4940 750 5040
rect 790 4940 890 5040
rect 930 4940 1030 5040
rect 1070 4940 1170 5040
rect 1210 4940 1310 5040
rect 2010 4940 2110 5040
rect 2150 4940 2250 5040
rect 2290 4940 2390 5040
rect 2430 4940 2530 5040
rect 2570 4940 2670 5040
rect 2710 4940 2810 5040
rect 2850 4940 2950 5040
rect 2990 4940 3090 5040
rect 3130 4940 3230 5040
rect 3270 4940 3370 5040
rect 3410 4940 3510 5040
rect -310 4150 -110 4650
rect -310 3610 -110 4110
rect 3430 4150 3630 4650
rect 3430 3610 3630 4110
<< ndiff >>
rect -30 7640 70 7650
rect -30 7620 0 7640
rect 40 7620 70 7640
rect -30 7610 70 7620
rect 140 7640 240 7650
rect 140 7620 170 7640
rect 210 7620 240 7640
rect 140 7610 240 7620
rect 310 7640 410 7650
rect 310 7620 340 7640
rect 380 7620 410 7640
rect 310 7610 410 7620
rect 480 7640 580 7650
rect 480 7620 510 7640
rect 550 7620 580 7640
rect 480 7610 580 7620
rect 650 7640 750 7650
rect 650 7620 680 7640
rect 720 7620 750 7640
rect 650 7610 750 7620
rect 820 7640 920 7650
rect 820 7620 850 7640
rect 890 7620 920 7640
rect 820 7610 920 7620
rect 990 7640 1090 7650
rect 990 7620 1020 7640
rect 1060 7620 1090 7640
rect 990 7610 1090 7620
rect 1160 7640 1260 7650
rect 1160 7620 1190 7640
rect 1230 7620 1260 7640
rect 1160 7610 1260 7620
rect 1330 7640 1430 7650
rect 1330 7620 1360 7640
rect 1400 7620 1430 7640
rect 1330 7610 1430 7620
rect 1500 7640 1600 7650
rect 1500 7620 1530 7640
rect 1570 7620 1600 7640
rect 1500 7610 1600 7620
rect 1720 7640 1820 7650
rect 1720 7620 1750 7640
rect 1790 7620 1820 7640
rect 1720 7610 1820 7620
rect 1890 7640 1990 7650
rect 1890 7620 1920 7640
rect 1960 7620 1990 7640
rect 1890 7610 1990 7620
rect 2060 7640 2160 7650
rect 2060 7620 2090 7640
rect 2130 7620 2160 7640
rect 2060 7610 2160 7620
rect 2230 7640 2330 7650
rect 2230 7620 2260 7640
rect 2300 7620 2330 7640
rect 2230 7610 2330 7620
rect 2400 7640 2500 7650
rect 2400 7620 2430 7640
rect 2470 7620 2500 7640
rect 2400 7610 2500 7620
rect 2570 7640 2670 7650
rect 2570 7620 2600 7640
rect 2640 7620 2670 7640
rect 2570 7610 2670 7620
rect 2740 7640 2840 7650
rect 2740 7620 2770 7640
rect 2810 7620 2840 7640
rect 2740 7610 2840 7620
rect 2910 7640 3010 7650
rect 2910 7620 2940 7640
rect 2980 7620 3010 7640
rect 2910 7610 3010 7620
rect 3080 7640 3180 7650
rect 3080 7620 3110 7640
rect 3150 7620 3180 7640
rect 3080 7610 3180 7620
rect 3250 7640 3350 7650
rect 3250 7620 3280 7640
rect 3320 7620 3350 7640
rect 3250 7610 3350 7620
rect -30 6600 70 6610
rect 140 6600 240 6610
rect 310 6600 410 6610
rect 480 6600 580 6610
rect 650 6600 750 6610
rect 820 6600 920 6610
rect 990 6600 1090 6610
rect 1160 6600 1260 6610
rect 1330 6600 1430 6610
rect 1500 6600 1600 6610
rect 1720 6600 1820 6610
rect 1890 6600 1990 6610
rect 2060 6600 2160 6610
rect 2230 6600 2330 6610
rect 2400 6600 2500 6610
rect 2570 6600 2670 6610
rect 2740 6600 2840 6610
rect 2910 6600 3010 6610
rect 3080 6600 3180 6610
rect 3250 6600 3350 6610
rect -30 6580 0 6600
rect 40 6580 170 6600
rect 210 6580 340 6600
rect 380 6580 510 6600
rect 550 6580 680 6600
rect 720 6580 850 6600
rect 890 6580 1020 6600
rect 1060 6580 1190 6600
rect 1230 6580 1360 6600
rect 1400 6580 1530 6600
rect 1570 6580 1750 6600
rect 1790 6580 1920 6600
rect 1960 6580 2090 6600
rect 2130 6580 2260 6600
rect 2300 6580 2430 6600
rect 2470 6580 2600 6600
rect 2640 6580 2770 6600
rect 2810 6580 2940 6600
rect 2980 6580 3110 6600
rect 3150 6580 3280 6600
rect 3320 6580 3350 6600
rect -30 6570 70 6580
rect 140 6570 240 6580
rect 310 6570 410 6580
rect 480 6570 580 6580
rect 650 6570 750 6580
rect 820 6570 920 6580
rect 990 6570 1090 6580
rect 1160 6570 1260 6580
rect 1330 6570 1430 6580
rect 1500 6570 1600 6580
rect 1720 6570 1820 6580
rect 1890 6570 1990 6580
rect 2060 6570 2160 6580
rect 2230 6570 2330 6580
rect 2400 6570 2500 6580
rect 2570 6570 2670 6580
rect 2740 6570 2840 6580
rect 2910 6570 3010 6580
rect 3080 6570 3180 6580
rect 3250 6570 3350 6580
rect -30 5560 70 5570
rect -30 5540 0 5560
rect 40 5540 70 5560
rect -30 5530 70 5540
rect -30 5490 -10 5530
rect 50 5490 70 5530
rect -30 5460 70 5490
rect 140 5560 240 5570
rect 140 5540 170 5560
rect 210 5540 240 5560
rect 140 5530 240 5540
rect 140 5490 160 5530
rect 220 5490 240 5530
rect 140 5460 240 5490
rect 310 5560 410 5570
rect 310 5540 340 5560
rect 380 5540 410 5560
rect 310 5530 410 5540
rect 310 5490 330 5530
rect 390 5490 410 5530
rect 310 5460 410 5490
rect 480 5560 580 5570
rect 480 5540 510 5560
rect 550 5540 580 5560
rect 480 5530 580 5540
rect 480 5490 500 5530
rect 560 5490 580 5530
rect 480 5460 580 5490
rect 650 5560 750 5570
rect 650 5540 680 5560
rect 720 5540 750 5560
rect 650 5530 750 5540
rect 650 5490 670 5530
rect 730 5490 750 5530
rect 650 5460 750 5490
rect 820 5560 920 5570
rect 820 5540 850 5560
rect 890 5540 920 5560
rect 820 5530 920 5540
rect 820 5490 840 5530
rect 900 5490 920 5530
rect 820 5460 920 5490
rect 990 5560 1090 5570
rect 990 5540 1020 5560
rect 1060 5540 1090 5560
rect 990 5530 1090 5540
rect 990 5490 1010 5530
rect 1070 5490 1090 5530
rect 990 5460 1090 5490
rect 1160 5560 1260 5570
rect 1160 5540 1190 5560
rect 1230 5540 1260 5560
rect 1160 5530 1260 5540
rect 1160 5490 1180 5530
rect 1240 5490 1260 5530
rect 1160 5460 1260 5490
rect 1330 5560 1430 5570
rect 1330 5540 1360 5560
rect 1400 5540 1430 5560
rect 1330 5530 1430 5540
rect 1330 5490 1350 5530
rect 1410 5490 1430 5530
rect 1330 5460 1430 5490
rect 1500 5560 1600 5570
rect 1500 5540 1530 5560
rect 1570 5540 1600 5560
rect 1500 5530 1600 5540
rect 1500 5490 1520 5530
rect 1580 5490 1600 5530
rect 1500 5460 1600 5490
rect 1720 5560 1820 5570
rect 1720 5540 1750 5560
rect 1790 5540 1820 5560
rect 1720 5530 1820 5540
rect 1720 5490 1740 5530
rect 1800 5490 1820 5530
rect 1720 5460 1820 5490
rect 1890 5560 1990 5570
rect 1890 5540 1920 5560
rect 1960 5540 1990 5560
rect 1890 5530 1990 5540
rect 1890 5490 1910 5530
rect 1970 5490 1990 5530
rect 1890 5460 1990 5490
rect 2060 5560 2160 5570
rect 2060 5540 2090 5560
rect 2130 5540 2160 5560
rect 2060 5530 2160 5540
rect 2060 5490 2080 5530
rect 2140 5490 2160 5530
rect 2060 5460 2160 5490
rect 2230 5560 2330 5570
rect 2230 5540 2260 5560
rect 2300 5540 2330 5560
rect 2230 5530 2330 5540
rect 2230 5490 2250 5530
rect 2310 5490 2330 5530
rect 2230 5460 2330 5490
rect 2400 5560 2500 5570
rect 2400 5540 2430 5560
rect 2470 5540 2500 5560
rect 2400 5530 2500 5540
rect 2400 5490 2420 5530
rect 2480 5490 2500 5530
rect 2400 5460 2500 5490
rect 2570 5560 2670 5570
rect 2570 5540 2600 5560
rect 2640 5540 2670 5560
rect 2570 5530 2670 5540
rect 2570 5490 2590 5530
rect 2650 5490 2670 5530
rect 2570 5460 2670 5490
rect 2740 5560 2840 5570
rect 2740 5540 2770 5560
rect 2810 5540 2840 5560
rect 2740 5530 2840 5540
rect 2740 5490 2760 5530
rect 2820 5490 2840 5530
rect 2740 5460 2840 5490
rect 2910 5560 3010 5570
rect 2910 5540 2940 5560
rect 2980 5540 3010 5560
rect 2910 5530 3010 5540
rect 2910 5490 2930 5530
rect 2990 5490 3010 5530
rect 2910 5460 3010 5490
rect 3080 5560 3180 5570
rect 3080 5540 3110 5560
rect 3150 5540 3180 5560
rect 3080 5530 3180 5540
rect 3080 5490 3100 5530
rect 3160 5490 3180 5530
rect 3080 5460 3180 5490
rect 3250 5560 3350 5570
rect 3250 5540 3280 5560
rect 3320 5540 3350 5560
rect 3250 5530 3350 5540
rect 3250 5490 3270 5530
rect 3330 5490 3350 5530
rect 3250 5460 3350 5490
rect -30 5350 70 5360
rect -30 5330 0 5350
rect 40 5330 70 5350
rect -30 5320 70 5330
rect 140 5350 240 5360
rect 140 5330 170 5350
rect 210 5330 240 5350
rect 140 5320 240 5330
rect 310 5350 410 5360
rect 310 5330 340 5350
rect 380 5330 410 5350
rect 310 5320 410 5330
rect 480 5350 580 5360
rect 480 5330 510 5350
rect 550 5330 580 5350
rect 480 5320 580 5330
rect 650 5350 750 5360
rect 650 5330 680 5350
rect 720 5330 750 5350
rect 650 5320 750 5330
rect 820 5350 920 5360
rect 820 5330 850 5350
rect 890 5330 920 5350
rect 820 5320 920 5330
rect 990 5350 1090 5360
rect 990 5330 1020 5350
rect 1060 5330 1090 5350
rect 990 5320 1090 5330
rect 1160 5350 1260 5360
rect 1160 5330 1190 5350
rect 1230 5330 1260 5350
rect 1160 5320 1260 5330
rect 1330 5350 1430 5360
rect 1330 5330 1360 5350
rect 1400 5330 1430 5350
rect 1330 5320 1430 5330
rect 1500 5350 1600 5360
rect 1500 5330 1530 5350
rect 1570 5330 1600 5350
rect 1500 5320 1600 5330
rect 1720 5350 1820 5360
rect 1720 5330 1750 5350
rect 1790 5330 1820 5350
rect 1720 5320 1820 5330
rect 1890 5350 1990 5360
rect 1890 5330 1920 5350
rect 1960 5330 1990 5350
rect 1890 5320 1990 5330
rect 2060 5350 2160 5360
rect 2060 5330 2090 5350
rect 2130 5330 2160 5350
rect 2060 5320 2160 5330
rect 2230 5350 2330 5360
rect 2230 5330 2260 5350
rect 2300 5330 2330 5350
rect 2230 5320 2330 5330
rect 2400 5350 2500 5360
rect 2400 5330 2430 5350
rect 2470 5330 2500 5350
rect 2400 5320 2500 5330
rect 2570 5350 2670 5360
rect 2570 5330 2600 5350
rect 2640 5330 2670 5350
rect 2570 5320 2670 5330
rect 2740 5350 2840 5360
rect 2740 5330 2770 5350
rect 2810 5330 2840 5350
rect 2740 5320 2840 5330
rect 2910 5350 3010 5360
rect 2910 5330 2940 5350
rect 2980 5330 3010 5350
rect 2910 5320 3010 5330
rect 3080 5350 3180 5360
rect 3080 5330 3110 5350
rect 3150 5330 3180 5350
rect 3080 5320 3180 5330
rect 3250 5350 3350 5360
rect 3250 5330 3280 5350
rect 3320 5330 3350 5350
rect 3250 5320 3350 5330
rect -30 4850 70 4860
rect -30 4830 0 4850
rect 40 4830 70 4850
rect -30 4820 70 4830
rect 140 4850 240 4860
rect 140 4830 170 4850
rect 210 4830 240 4850
rect 140 4820 240 4830
rect 310 4850 410 4860
rect 310 4830 340 4850
rect 380 4830 410 4850
rect 310 4820 410 4830
rect 480 4850 580 4860
rect 480 4830 510 4850
rect 550 4830 580 4850
rect 480 4820 580 4830
rect 650 4850 750 4860
rect 650 4830 680 4850
rect 720 4830 750 4850
rect 650 4820 750 4830
rect 820 4850 920 4860
rect 820 4830 850 4850
rect 890 4830 920 4850
rect 820 4820 920 4830
rect 990 4850 1090 4860
rect 990 4830 1020 4850
rect 1060 4830 1090 4850
rect 990 4820 1090 4830
rect 1160 4850 1260 4860
rect 1160 4830 1190 4850
rect 1230 4830 1260 4850
rect 1160 4820 1260 4830
rect 1330 4850 1430 4860
rect 1330 4830 1360 4850
rect 1400 4830 1430 4850
rect 1330 4820 1430 4830
rect 1500 4850 1600 4860
rect 1500 4830 1530 4850
rect 1570 4830 1600 4850
rect 1500 4820 1600 4830
rect 1720 4850 1820 4860
rect 1720 4830 1750 4850
rect 1790 4830 1820 4850
rect 1720 4820 1820 4830
rect 1890 4850 1990 4860
rect 1890 4830 1920 4850
rect 1960 4830 1990 4850
rect 1890 4820 1990 4830
rect 2060 4850 2160 4860
rect 2060 4830 2090 4850
rect 2130 4830 2160 4850
rect 2060 4820 2160 4830
rect 2230 4850 2330 4860
rect 2230 4830 2260 4850
rect 2300 4830 2330 4850
rect 2230 4820 2330 4830
rect 2400 4850 2500 4860
rect 2400 4830 2430 4850
rect 2470 4830 2500 4850
rect 2400 4820 2500 4830
rect 2570 4850 2670 4860
rect 2570 4830 2600 4850
rect 2640 4830 2670 4850
rect 2570 4820 2670 4830
rect 2740 4850 2840 4860
rect 2740 4830 2770 4850
rect 2810 4830 2840 4850
rect 2740 4820 2840 4830
rect 2910 4850 3010 4860
rect 2910 4830 2940 4850
rect 2980 4830 3010 4850
rect 2910 4820 3010 4830
rect 3080 4850 3180 4860
rect 3080 4830 3110 4850
rect 3150 4830 3180 4850
rect 3080 4820 3180 4830
rect 3250 4850 3350 4860
rect 3250 4830 3280 4850
rect 3320 4830 3350 4850
rect 3250 4820 3350 4830
rect -30 4690 70 4720
rect -30 4650 -10 4690
rect 50 4650 70 4690
rect -30 4640 70 4650
rect -30 4620 0 4640
rect 40 4620 70 4640
rect -30 4610 70 4620
rect 140 4690 240 4720
rect 140 4650 160 4690
rect 220 4650 240 4690
rect 140 4640 240 4650
rect 140 4620 170 4640
rect 210 4620 240 4640
rect 140 4610 240 4620
rect 310 4690 410 4720
rect 310 4650 330 4690
rect 390 4650 410 4690
rect 310 4640 410 4650
rect 310 4620 340 4640
rect 380 4620 410 4640
rect 310 4610 410 4620
rect 480 4690 580 4720
rect 480 4650 500 4690
rect 560 4650 580 4690
rect 480 4640 580 4650
rect 480 4620 510 4640
rect 550 4620 580 4640
rect 480 4610 580 4620
rect 650 4690 750 4720
rect 650 4650 670 4690
rect 730 4650 750 4690
rect 650 4640 750 4650
rect 650 4620 680 4640
rect 720 4620 750 4640
rect 650 4610 750 4620
rect 820 4690 920 4720
rect 820 4650 840 4690
rect 900 4650 920 4690
rect 820 4640 920 4650
rect 820 4620 850 4640
rect 890 4620 920 4640
rect 820 4610 920 4620
rect 990 4690 1090 4720
rect 990 4650 1010 4690
rect 1070 4650 1090 4690
rect 990 4640 1090 4650
rect 990 4620 1020 4640
rect 1060 4620 1090 4640
rect 990 4610 1090 4620
rect 1160 4690 1260 4720
rect 1160 4650 1180 4690
rect 1240 4650 1260 4690
rect 1160 4640 1260 4650
rect 1160 4620 1190 4640
rect 1230 4620 1260 4640
rect 1160 4610 1260 4620
rect 1330 4690 1430 4720
rect 1330 4650 1350 4690
rect 1410 4650 1430 4690
rect 1330 4640 1430 4650
rect 1330 4620 1360 4640
rect 1400 4620 1430 4640
rect 1330 4610 1430 4620
rect 1500 4690 1600 4720
rect 1500 4650 1520 4690
rect 1580 4650 1600 4690
rect 1500 4640 1600 4650
rect 1500 4620 1530 4640
rect 1570 4620 1600 4640
rect 1500 4610 1600 4620
rect 1720 4690 1820 4720
rect 1720 4650 1740 4690
rect 1800 4650 1820 4690
rect 1720 4640 1820 4650
rect 1720 4620 1750 4640
rect 1790 4620 1820 4640
rect 1720 4610 1820 4620
rect 1890 4690 1990 4720
rect 1890 4650 1910 4690
rect 1970 4650 1990 4690
rect 1890 4640 1990 4650
rect 1890 4620 1920 4640
rect 1960 4620 1990 4640
rect 1890 4610 1990 4620
rect 2060 4690 2160 4720
rect 2060 4650 2080 4690
rect 2140 4650 2160 4690
rect 2060 4640 2160 4650
rect 2060 4620 2090 4640
rect 2130 4620 2160 4640
rect 2060 4610 2160 4620
rect 2230 4690 2330 4720
rect 2230 4650 2250 4690
rect 2310 4650 2330 4690
rect 2230 4640 2330 4650
rect 2230 4620 2260 4640
rect 2300 4620 2330 4640
rect 2230 4610 2330 4620
rect 2400 4690 2500 4720
rect 2400 4650 2420 4690
rect 2480 4650 2500 4690
rect 2400 4640 2500 4650
rect 2400 4620 2430 4640
rect 2470 4620 2500 4640
rect 2400 4610 2500 4620
rect 2570 4690 2670 4720
rect 2570 4650 2590 4690
rect 2650 4650 2670 4690
rect 2570 4640 2670 4650
rect 2570 4620 2600 4640
rect 2640 4620 2670 4640
rect 2570 4610 2670 4620
rect 2740 4690 2840 4720
rect 2740 4650 2760 4690
rect 2820 4650 2840 4690
rect 2740 4640 2840 4650
rect 2740 4620 2770 4640
rect 2810 4620 2840 4640
rect 2740 4610 2840 4620
rect 2910 4690 3010 4720
rect 2910 4650 2930 4690
rect 2990 4650 3010 4690
rect 2910 4640 3010 4650
rect 2910 4620 2940 4640
rect 2980 4620 3010 4640
rect 2910 4610 3010 4620
rect 3080 4690 3180 4720
rect 3080 4650 3100 4690
rect 3160 4650 3180 4690
rect 3080 4640 3180 4650
rect 3080 4620 3110 4640
rect 3150 4620 3180 4640
rect 3080 4610 3180 4620
rect 3250 4690 3350 4720
rect 3250 4650 3270 4690
rect 3330 4650 3350 4690
rect 3250 4640 3350 4650
rect 3250 4620 3280 4640
rect 3320 4620 3350 4640
rect 3250 4610 3350 4620
rect -30 3600 70 3610
rect 140 3600 240 3610
rect 310 3600 410 3610
rect 480 3600 580 3610
rect 650 3600 750 3610
rect 820 3600 920 3610
rect 990 3600 1090 3610
rect 1160 3600 1260 3610
rect 1330 3600 1430 3610
rect 1500 3600 1600 3610
rect 1720 3600 1820 3610
rect 1890 3600 1990 3610
rect 2060 3600 2160 3610
rect 2230 3600 2330 3610
rect 2400 3600 2500 3610
rect 2570 3600 2670 3610
rect 2740 3600 2840 3610
rect 2910 3600 3010 3610
rect 3080 3600 3180 3610
rect 3250 3600 3350 3610
rect -30 3580 0 3600
rect 40 3580 170 3600
rect 210 3580 340 3600
rect 380 3580 510 3600
rect 550 3580 680 3600
rect 720 3580 850 3600
rect 890 3580 1020 3600
rect 1060 3580 1190 3600
rect 1230 3580 1360 3600
rect 1400 3580 1530 3600
rect 1570 3580 1750 3600
rect 1790 3580 1920 3600
rect 1960 3580 2090 3600
rect 2130 3580 2260 3600
rect 2300 3580 2430 3600
rect 2470 3580 2600 3600
rect 2640 3580 2770 3600
rect 2810 3580 2940 3600
rect 2980 3580 3110 3600
rect 3150 3580 3280 3600
rect 3320 3580 3350 3600
rect -30 3570 70 3580
rect 140 3570 240 3580
rect 310 3570 410 3580
rect 480 3570 580 3580
rect 650 3570 750 3580
rect 820 3570 920 3580
rect 990 3570 1090 3580
rect 1160 3570 1260 3580
rect 1330 3570 1430 3580
rect 1500 3570 1600 3580
rect 1720 3570 1820 3580
rect 1890 3570 1990 3580
rect 2060 3570 2160 3580
rect 2230 3570 2330 3580
rect 2400 3570 2500 3580
rect 2570 3570 2670 3580
rect 2740 3570 2840 3580
rect 2910 3570 3010 3580
rect 3080 3570 3180 3580
rect 3250 3570 3350 3580
rect -30 2560 70 2570
rect -30 2540 0 2560
rect 40 2540 70 2560
rect -30 2530 70 2540
rect 140 2560 240 2570
rect 140 2540 170 2560
rect 210 2540 240 2560
rect 140 2530 240 2540
rect 310 2560 410 2570
rect 310 2540 340 2560
rect 380 2540 410 2560
rect 310 2530 410 2540
rect 480 2560 580 2570
rect 480 2540 510 2560
rect 550 2540 580 2560
rect 480 2530 580 2540
rect 650 2560 750 2570
rect 650 2540 680 2560
rect 720 2540 750 2560
rect 650 2530 750 2540
rect 820 2560 920 2570
rect 820 2540 850 2560
rect 890 2540 920 2560
rect 820 2530 920 2540
rect 990 2560 1090 2570
rect 990 2540 1020 2560
rect 1060 2540 1090 2560
rect 990 2530 1090 2540
rect 1160 2560 1260 2570
rect 1160 2540 1190 2560
rect 1230 2540 1260 2560
rect 1160 2530 1260 2540
rect 1330 2560 1430 2570
rect 1330 2540 1360 2560
rect 1400 2540 1430 2560
rect 1330 2530 1430 2540
rect 1500 2560 1600 2570
rect 1500 2540 1530 2560
rect 1570 2540 1600 2560
rect 1500 2530 1600 2540
rect 1720 2560 1820 2570
rect 1720 2540 1750 2560
rect 1790 2540 1820 2560
rect 1720 2530 1820 2540
rect 1890 2560 1990 2570
rect 1890 2540 1920 2560
rect 1960 2540 1990 2560
rect 1890 2530 1990 2540
rect 2060 2560 2160 2570
rect 2060 2540 2090 2560
rect 2130 2540 2160 2560
rect 2060 2530 2160 2540
rect 2230 2560 2330 2570
rect 2230 2540 2260 2560
rect 2300 2540 2330 2560
rect 2230 2530 2330 2540
rect 2400 2560 2500 2570
rect 2400 2540 2430 2560
rect 2470 2540 2500 2560
rect 2400 2530 2500 2540
rect 2570 2560 2670 2570
rect 2570 2540 2600 2560
rect 2640 2540 2670 2560
rect 2570 2530 2670 2540
rect 2740 2560 2840 2570
rect 2740 2540 2770 2560
rect 2810 2540 2840 2560
rect 2740 2530 2840 2540
rect 2910 2560 3010 2570
rect 2910 2540 2940 2560
rect 2980 2540 3010 2560
rect 2910 2530 3010 2540
rect 3080 2560 3180 2570
rect 3080 2540 3110 2560
rect 3150 2540 3180 2560
rect 3080 2530 3180 2540
rect 3250 2560 3350 2570
rect 3250 2540 3280 2560
rect 3320 2540 3350 2560
rect 3250 2530 3350 2540
<< pdiff >>
rect -310 6600 -110 6610
rect -310 6580 -230 6600
rect -190 6580 -110 6600
rect -310 6570 -110 6580
rect 3430 6600 3630 6610
rect 3430 6580 3510 6600
rect 3550 6580 3630 6600
rect 3430 6570 3630 6580
rect -310 6060 -110 6070
rect -310 6040 -230 6060
rect -190 6040 -110 6060
rect -310 6030 -110 6040
rect -310 5520 -110 5530
rect -310 5500 -230 5520
rect -190 5500 -110 5520
rect -310 5490 -110 5500
rect 3430 6060 3630 6070
rect 3430 6040 3510 6060
rect 3550 6040 3630 6060
rect 3430 6030 3630 6040
rect 3430 5520 3630 5530
rect 3430 5500 3510 5520
rect 3550 5500 3630 5520
rect 3430 5490 3630 5500
rect 1520 5240 1560 5250
rect 1760 5240 1800 5250
rect -270 5220 -190 5240
rect -230 5210 -190 5220
rect -230 5170 -220 5210
rect -200 5170 -190 5210
rect -230 5160 -190 5170
rect -270 5140 -190 5160
rect -90 5210 -50 5240
rect -90 5170 -80 5210
rect -60 5170 -50 5210
rect -90 5140 -50 5170
rect 50 5210 90 5240
rect 50 5170 60 5210
rect 80 5170 90 5210
rect 50 5140 90 5170
rect 190 5210 230 5240
rect 190 5170 200 5210
rect 220 5170 230 5210
rect 190 5140 230 5170
rect 330 5210 370 5240
rect 330 5170 340 5210
rect 360 5170 370 5210
rect 330 5140 370 5170
rect 470 5210 510 5240
rect 470 5170 480 5210
rect 500 5170 510 5210
rect 470 5140 510 5170
rect 610 5210 650 5240
rect 610 5170 620 5210
rect 640 5170 650 5210
rect 610 5140 650 5170
rect 750 5210 790 5240
rect 750 5170 760 5210
rect 780 5170 790 5210
rect 750 5140 790 5170
rect 890 5210 930 5240
rect 890 5170 900 5210
rect 920 5170 930 5210
rect 890 5140 930 5170
rect 1030 5210 1070 5240
rect 1030 5170 1040 5210
rect 1060 5170 1070 5210
rect 1030 5140 1070 5170
rect 1170 5210 1210 5240
rect 1170 5170 1180 5210
rect 1200 5170 1210 5210
rect 1170 5140 1210 5170
rect 1310 5210 1350 5240
rect 1520 5220 1530 5240
rect 1550 5220 1770 5240
rect 1790 5220 1800 5240
rect 1520 5210 1800 5220
rect 1970 5210 2010 5240
rect 1310 5170 1320 5210
rect 1340 5170 1350 5210
rect 1310 5140 1350 5170
rect 1520 5170 1800 5180
rect 1520 5150 1530 5170
rect 1550 5150 1770 5170
rect 1790 5150 1800 5170
rect 1520 5140 1800 5150
rect 1970 5170 1980 5210
rect 2000 5170 2010 5210
rect 1970 5140 2010 5170
rect 2110 5210 2150 5240
rect 2110 5170 2120 5210
rect 2140 5170 2150 5210
rect 2110 5140 2150 5170
rect 2250 5210 2290 5240
rect 2250 5170 2260 5210
rect 2280 5170 2290 5210
rect 2250 5140 2290 5170
rect 2390 5210 2430 5240
rect 2390 5170 2400 5210
rect 2420 5170 2430 5210
rect 2390 5140 2430 5170
rect 2530 5210 2570 5240
rect 2530 5170 2540 5210
rect 2560 5170 2570 5210
rect 2530 5140 2570 5170
rect 2670 5210 2710 5240
rect 2670 5170 2680 5210
rect 2700 5170 2710 5210
rect 2670 5140 2710 5170
rect 2810 5210 2850 5240
rect 2810 5170 2820 5210
rect 2840 5170 2850 5210
rect 2810 5140 2850 5170
rect 2950 5210 2990 5240
rect 2950 5170 2960 5210
rect 2980 5170 2990 5210
rect 2950 5140 2990 5170
rect 3090 5210 3130 5240
rect 3090 5170 3100 5210
rect 3120 5170 3130 5210
rect 3090 5140 3130 5170
rect 3230 5210 3270 5240
rect 3230 5170 3240 5210
rect 3260 5170 3270 5210
rect 3230 5140 3270 5170
rect 3370 5210 3410 5240
rect 3370 5170 3380 5210
rect 3400 5170 3410 5210
rect 3370 5140 3410 5170
rect 3510 5220 3590 5240
rect 3510 5210 3550 5220
rect 3510 5170 3520 5210
rect 3540 5170 3550 5210
rect 3510 5160 3550 5170
rect 3510 5140 3590 5160
rect 1180 5040 1200 5140
rect 1320 5040 1340 5140
rect 1520 5100 1800 5110
rect 1520 5080 1530 5100
rect 1550 5080 1770 5100
rect 1790 5080 1800 5100
rect 1520 5070 1800 5080
rect 1980 5040 2000 5140
rect 2120 5040 2140 5140
rect -270 5020 -190 5040
rect -230 5010 -190 5020
rect -230 4970 -220 5010
rect -200 4970 -190 5010
rect -230 4960 -190 4970
rect -270 4940 -190 4960
rect -90 5010 -50 5040
rect -90 4970 -80 5010
rect -60 4970 -50 5010
rect -90 4940 -50 4970
rect 50 5010 90 5040
rect 50 4970 60 5010
rect 80 4970 90 5010
rect 50 4940 90 4970
rect 190 5010 230 5040
rect 190 4970 200 5010
rect 220 4970 230 5010
rect 190 4940 230 4970
rect 330 5010 370 5040
rect 330 4970 340 5010
rect 360 4970 370 5010
rect 330 4940 370 4970
rect 470 5010 510 5040
rect 470 4970 480 5010
rect 500 4970 510 5010
rect 470 4940 510 4970
rect 610 5010 650 5040
rect 610 4970 620 5010
rect 640 4970 650 5010
rect 610 4940 650 4970
rect 750 5010 790 5040
rect 750 4970 760 5010
rect 780 4970 790 5010
rect 750 4940 790 4970
rect 890 5010 930 5040
rect 890 4970 900 5010
rect 920 4970 930 5010
rect 890 4940 930 4970
rect 1030 5010 1070 5040
rect 1030 4970 1040 5010
rect 1060 4970 1070 5010
rect 1030 4940 1070 4970
rect 1170 5010 1210 5040
rect 1170 4970 1180 5010
rect 1200 4970 1210 5010
rect 1170 4940 1210 4970
rect 1310 5010 1350 5040
rect 1310 4970 1320 5010
rect 1340 4970 1350 5010
rect 1520 5030 1800 5040
rect 1520 5010 1530 5030
rect 1550 5010 1770 5030
rect 1790 5010 1800 5030
rect 1520 5000 1800 5010
rect 1970 5010 2010 5040
rect 1970 4970 1980 5010
rect 2000 4970 2010 5010
rect 1310 4940 1350 4970
rect 1520 4960 1800 4970
rect 1520 4940 1530 4960
rect 1550 4940 1770 4960
rect 1790 4940 1800 4960
rect 1970 4940 2010 4970
rect 2110 5010 2150 5040
rect 2110 4970 2120 5010
rect 2140 4970 2150 5010
rect 2110 4940 2150 4970
rect 2250 5010 2290 5040
rect 2250 4970 2260 5010
rect 2280 4970 2290 5010
rect 2250 4940 2290 4970
rect 2390 5010 2430 5040
rect 2390 4970 2400 5010
rect 2420 4970 2430 5010
rect 2390 4940 2430 4970
rect 2530 5010 2570 5040
rect 2530 4970 2540 5010
rect 2560 4970 2570 5010
rect 2530 4940 2570 4970
rect 2670 5010 2710 5040
rect 2670 4970 2680 5010
rect 2700 4970 2710 5010
rect 2670 4940 2710 4970
rect 2810 5010 2850 5040
rect 2810 4970 2820 5010
rect 2840 4970 2850 5010
rect 2810 4940 2850 4970
rect 2950 5010 2990 5040
rect 2950 4970 2960 5010
rect 2980 4970 2990 5010
rect 2950 4940 2990 4970
rect 3090 5010 3130 5040
rect 3090 4970 3100 5010
rect 3120 4970 3130 5010
rect 3090 4940 3130 4970
rect 3230 5010 3270 5040
rect 3230 4970 3240 5010
rect 3260 4970 3270 5010
rect 3230 4940 3270 4970
rect 3370 5010 3410 5040
rect 3370 4970 3380 5010
rect 3400 4970 3410 5010
rect 3370 4940 3410 4970
rect 3510 5020 3590 5040
rect 3510 5010 3550 5020
rect 3510 4970 3520 5010
rect 3540 4970 3550 5010
rect 3510 4960 3550 4970
rect 3510 4940 3590 4960
rect 1520 4930 1560 4940
rect 1760 4930 1800 4940
rect -310 4680 -110 4690
rect -310 4660 -230 4680
rect -190 4660 -110 4680
rect -310 4650 -110 4660
rect -310 4140 -110 4150
rect -310 4120 -230 4140
rect -190 4120 -110 4140
rect -310 4110 -110 4120
rect 3430 4680 3630 4690
rect 3430 4660 3510 4680
rect 3550 4660 3630 4680
rect 3430 4650 3630 4660
rect 3430 4140 3630 4150
rect 3430 4120 3510 4140
rect 3550 4120 3630 4140
rect 3430 4110 3630 4120
rect -310 3600 -110 3610
rect -310 3580 -230 3600
rect -190 3580 -110 3600
rect -310 3570 -110 3580
rect 3430 3600 3630 3610
rect 3430 3580 3510 3600
rect 3550 3580 3630 3600
rect 3430 3570 3630 3580
<< ndiffc >>
rect 0 7620 40 7640
rect 170 7620 210 7640
rect 340 7620 380 7640
rect 510 7620 550 7640
rect 680 7620 720 7640
rect 850 7620 890 7640
rect 1020 7620 1060 7640
rect 1190 7620 1230 7640
rect 1360 7620 1400 7640
rect 1530 7620 1570 7640
rect 1750 7620 1790 7640
rect 1920 7620 1960 7640
rect 2090 7620 2130 7640
rect 2260 7620 2300 7640
rect 2430 7620 2470 7640
rect 2600 7620 2640 7640
rect 2770 7620 2810 7640
rect 2940 7620 2980 7640
rect 3110 7620 3150 7640
rect 3280 7620 3320 7640
rect 0 6580 40 6600
rect 170 6580 210 6600
rect 340 6580 380 6600
rect 510 6580 550 6600
rect 680 6580 720 6600
rect 850 6580 890 6600
rect 1020 6580 1060 6600
rect 1190 6580 1230 6600
rect 1360 6580 1400 6600
rect 1530 6580 1570 6600
rect 1750 6580 1790 6600
rect 1920 6580 1960 6600
rect 2090 6580 2130 6600
rect 2260 6580 2300 6600
rect 2430 6580 2470 6600
rect 2600 6580 2640 6600
rect 2770 6580 2810 6600
rect 2940 6580 2980 6600
rect 3110 6580 3150 6600
rect 3280 6580 3320 6600
rect 0 5540 40 5560
rect 170 5540 210 5560
rect 340 5540 380 5560
rect 510 5540 550 5560
rect 680 5540 720 5560
rect 850 5540 890 5560
rect 1020 5540 1060 5560
rect 1190 5540 1230 5560
rect 1360 5540 1400 5560
rect 1530 5540 1570 5560
rect 1750 5540 1790 5560
rect 1920 5540 1960 5560
rect 2090 5540 2130 5560
rect 2260 5540 2300 5560
rect 2430 5540 2470 5560
rect 2600 5540 2640 5560
rect 2770 5540 2810 5560
rect 2940 5540 2980 5560
rect 3110 5540 3150 5560
rect 3280 5540 3320 5560
rect 0 5330 40 5350
rect 170 5330 210 5350
rect 340 5330 380 5350
rect 510 5330 550 5350
rect 680 5330 720 5350
rect 850 5330 890 5350
rect 1020 5330 1060 5350
rect 1190 5330 1230 5350
rect 1360 5330 1400 5350
rect 1530 5330 1570 5350
rect 1750 5330 1790 5350
rect 1920 5330 1960 5350
rect 2090 5330 2130 5350
rect 2260 5330 2300 5350
rect 2430 5330 2470 5350
rect 2600 5330 2640 5350
rect 2770 5330 2810 5350
rect 2940 5330 2980 5350
rect 3110 5330 3150 5350
rect 3280 5330 3320 5350
rect 0 4830 40 4850
rect 170 4830 210 4850
rect 340 4830 380 4850
rect 510 4830 550 4850
rect 680 4830 720 4850
rect 850 4830 890 4850
rect 1020 4830 1060 4850
rect 1190 4830 1230 4850
rect 1360 4830 1400 4850
rect 1530 4830 1570 4850
rect 1750 4830 1790 4850
rect 1920 4830 1960 4850
rect 2090 4830 2130 4850
rect 2260 4830 2300 4850
rect 2430 4830 2470 4850
rect 2600 4830 2640 4850
rect 2770 4830 2810 4850
rect 2940 4830 2980 4850
rect 3110 4830 3150 4850
rect 3280 4830 3320 4850
rect 0 4620 40 4640
rect 170 4620 210 4640
rect 340 4620 380 4640
rect 510 4620 550 4640
rect 680 4620 720 4640
rect 850 4620 890 4640
rect 1020 4620 1060 4640
rect 1190 4620 1230 4640
rect 1360 4620 1400 4640
rect 1530 4620 1570 4640
rect 1750 4620 1790 4640
rect 1920 4620 1960 4640
rect 2090 4620 2130 4640
rect 2260 4620 2300 4640
rect 2430 4620 2470 4640
rect 2600 4620 2640 4640
rect 2770 4620 2810 4640
rect 2940 4620 2980 4640
rect 3110 4620 3150 4640
rect 3280 4620 3320 4640
rect 0 3580 40 3600
rect 170 3580 210 3600
rect 340 3580 380 3600
rect 510 3580 550 3600
rect 680 3580 720 3600
rect 850 3580 890 3600
rect 1020 3580 1060 3600
rect 1190 3580 1230 3600
rect 1360 3580 1400 3600
rect 1530 3580 1570 3600
rect 1750 3580 1790 3600
rect 1920 3580 1960 3600
rect 2090 3580 2130 3600
rect 2260 3580 2300 3600
rect 2430 3580 2470 3600
rect 2600 3580 2640 3600
rect 2770 3580 2810 3600
rect 2940 3580 2980 3600
rect 3110 3580 3150 3600
rect 3280 3580 3320 3600
rect 0 2540 40 2560
rect 170 2540 210 2560
rect 340 2540 380 2560
rect 510 2540 550 2560
rect 680 2540 720 2560
rect 850 2540 890 2560
rect 1020 2540 1060 2560
rect 1190 2540 1230 2560
rect 1360 2540 1400 2560
rect 1530 2540 1570 2560
rect 1750 2540 1790 2560
rect 1920 2540 1960 2560
rect 2090 2540 2130 2560
rect 2260 2540 2300 2560
rect 2430 2540 2470 2560
rect 2600 2540 2640 2560
rect 2770 2540 2810 2560
rect 2940 2540 2980 2560
rect 3110 2540 3150 2560
rect 3280 2540 3320 2560
<< pdiffc >>
rect -230 6580 -190 6600
rect 3510 6580 3550 6600
rect -230 6040 -190 6060
rect -230 5500 -190 5520
rect 3510 6040 3550 6060
rect 3510 5500 3550 5520
rect -220 5170 -200 5210
rect -80 5170 -60 5210
rect 60 5170 80 5210
rect 200 5170 220 5210
rect 340 5170 360 5210
rect 480 5170 500 5210
rect 620 5170 640 5210
rect 760 5170 780 5210
rect 900 5170 920 5210
rect 1040 5170 1060 5210
rect 1180 5170 1200 5210
rect 1530 5220 1550 5240
rect 1770 5220 1790 5240
rect 1320 5170 1340 5210
rect 1530 5150 1550 5170
rect 1770 5150 1790 5170
rect 1980 5170 2000 5210
rect 2120 5170 2140 5210
rect 2260 5170 2280 5210
rect 2400 5170 2420 5210
rect 2540 5170 2560 5210
rect 2680 5170 2700 5210
rect 2820 5170 2840 5210
rect 2960 5170 2980 5210
rect 3100 5170 3120 5210
rect 3240 5170 3260 5210
rect 3380 5170 3400 5210
rect 3520 5170 3540 5210
rect 1530 5080 1550 5100
rect 1770 5080 1790 5100
rect -220 4970 -200 5010
rect -80 4970 -60 5010
rect 60 4970 80 5010
rect 200 4970 220 5010
rect 340 4970 360 5010
rect 480 4970 500 5010
rect 620 4970 640 5010
rect 760 4970 780 5010
rect 900 4970 920 5010
rect 1040 4970 1060 5010
rect 1180 4970 1200 5010
rect 1320 4970 1340 5010
rect 1530 5010 1550 5030
rect 1770 5010 1790 5030
rect 1980 4970 2000 5010
rect 1530 4940 1550 4960
rect 1770 4940 1790 4960
rect 2120 4970 2140 5010
rect 2260 4970 2280 5010
rect 2400 4970 2420 5010
rect 2540 4970 2560 5010
rect 2680 4970 2700 5010
rect 2820 4970 2840 5010
rect 2960 4970 2980 5010
rect 3100 4970 3120 5010
rect 3240 4970 3260 5010
rect 3380 4970 3400 5010
rect 3520 4970 3540 5010
rect -230 4660 -190 4680
rect -230 4120 -190 4140
rect 3510 4660 3550 4680
rect 3510 4120 3550 4140
rect -230 3580 -190 3600
rect 3510 3580 3550 3600
<< psubdiff >>
rect -30 7660 0 7680
rect 40 7660 70 7680
rect -30 7650 70 7660
rect 140 7660 170 7680
rect 210 7660 240 7680
rect 140 7650 240 7660
rect 310 7660 340 7680
rect 380 7660 410 7680
rect 310 7650 410 7660
rect 480 7660 510 7680
rect 550 7660 580 7680
rect 480 7650 580 7660
rect 650 7660 680 7680
rect 720 7660 750 7680
rect 650 7650 750 7660
rect 820 7660 850 7680
rect 890 7660 920 7680
rect 820 7650 920 7660
rect 990 7660 1020 7680
rect 1060 7660 1090 7680
rect 990 7650 1090 7660
rect 1160 7660 1190 7680
rect 1230 7660 1260 7680
rect 1160 7650 1260 7660
rect 1330 7660 1360 7680
rect 1400 7660 1430 7680
rect 1330 7650 1430 7660
rect 1500 7660 1530 7680
rect 1570 7660 1600 7680
rect 1500 7650 1600 7660
rect 1720 7660 1750 7680
rect 1790 7660 1820 7680
rect 1720 7650 1820 7660
rect 1890 7660 1920 7680
rect 1960 7660 1990 7680
rect 1890 7650 1990 7660
rect 2060 7660 2090 7680
rect 2130 7660 2160 7680
rect 2060 7650 2160 7660
rect 2230 7660 2260 7680
rect 2300 7660 2330 7680
rect 2230 7650 2330 7660
rect 2400 7660 2430 7680
rect 2470 7660 2500 7680
rect 2400 7650 2500 7660
rect 2570 7660 2600 7680
rect 2640 7660 2670 7680
rect 2570 7650 2670 7660
rect 2740 7660 2770 7680
rect 2810 7660 2840 7680
rect 2740 7650 2840 7660
rect 2910 7660 2940 7680
rect 2980 7660 3010 7680
rect 2910 7650 3010 7660
rect 3080 7660 3110 7680
rect 3150 7660 3180 7680
rect 3080 7650 3180 7660
rect 3250 7660 3280 7680
rect 3320 7660 3350 7680
rect 3250 7650 3350 7660
rect -10 5520 50 5530
rect -10 5500 0 5520
rect 40 5500 50 5520
rect -10 5490 50 5500
rect 160 5520 220 5530
rect 160 5500 170 5520
rect 210 5500 220 5520
rect 160 5490 220 5500
rect 330 5520 390 5530
rect 330 5500 340 5520
rect 380 5500 390 5520
rect 330 5490 390 5500
rect 500 5520 560 5530
rect 500 5500 510 5520
rect 550 5500 560 5520
rect 500 5490 560 5500
rect 670 5520 730 5530
rect 670 5500 680 5520
rect 720 5500 730 5520
rect 670 5490 730 5500
rect 840 5520 900 5530
rect 840 5500 850 5520
rect 890 5500 900 5520
rect 840 5490 900 5500
rect 1010 5520 1070 5530
rect 1010 5500 1020 5520
rect 1060 5500 1070 5520
rect 1010 5490 1070 5500
rect 1180 5520 1240 5530
rect 1180 5500 1190 5520
rect 1230 5500 1240 5520
rect 1180 5490 1240 5500
rect 1350 5520 1410 5530
rect 1350 5500 1360 5520
rect 1400 5500 1410 5520
rect 1350 5490 1410 5500
rect 1520 5520 1580 5530
rect 1520 5500 1530 5520
rect 1570 5500 1580 5520
rect 1520 5490 1580 5500
rect 1740 5520 1800 5530
rect 1740 5500 1750 5520
rect 1790 5500 1800 5520
rect 1740 5490 1800 5500
rect 1910 5520 1970 5530
rect 1910 5500 1920 5520
rect 1960 5500 1970 5520
rect 1910 5490 1970 5500
rect 2080 5520 2140 5530
rect 2080 5500 2090 5520
rect 2130 5500 2140 5520
rect 2080 5490 2140 5500
rect 2250 5520 2310 5530
rect 2250 5500 2260 5520
rect 2300 5500 2310 5520
rect 2250 5490 2310 5500
rect 2420 5520 2480 5530
rect 2420 5500 2430 5520
rect 2470 5500 2480 5520
rect 2420 5490 2480 5500
rect 2590 5520 2650 5530
rect 2590 5500 2600 5520
rect 2640 5500 2650 5520
rect 2590 5490 2650 5500
rect 2760 5520 2820 5530
rect 2760 5500 2770 5520
rect 2810 5500 2820 5520
rect 2760 5490 2820 5500
rect 2930 5520 2990 5530
rect 2930 5500 2940 5520
rect 2980 5500 2990 5520
rect 2930 5490 2990 5500
rect 3100 5520 3160 5530
rect 3100 5500 3110 5520
rect 3150 5500 3160 5520
rect 3100 5490 3160 5500
rect 3270 5520 3330 5530
rect 3270 5500 3280 5520
rect 3320 5500 3330 5520
rect 3270 5490 3330 5500
rect -10 4680 50 4690
rect -10 4660 0 4680
rect 40 4660 50 4680
rect -10 4650 50 4660
rect 160 4680 220 4690
rect 160 4660 170 4680
rect 210 4660 220 4680
rect 160 4650 220 4660
rect 330 4680 390 4690
rect 330 4660 340 4680
rect 380 4660 390 4680
rect 330 4650 390 4660
rect 500 4680 560 4690
rect 500 4660 510 4680
rect 550 4660 560 4680
rect 500 4650 560 4660
rect 670 4680 730 4690
rect 670 4660 680 4680
rect 720 4660 730 4680
rect 670 4650 730 4660
rect 840 4680 900 4690
rect 840 4660 850 4680
rect 890 4660 900 4680
rect 840 4650 900 4660
rect 1010 4680 1070 4690
rect 1010 4660 1020 4680
rect 1060 4660 1070 4680
rect 1010 4650 1070 4660
rect 1180 4680 1240 4690
rect 1180 4660 1190 4680
rect 1230 4660 1240 4680
rect 1180 4650 1240 4660
rect 1350 4680 1410 4690
rect 1350 4660 1360 4680
rect 1400 4660 1410 4680
rect 1350 4650 1410 4660
rect 1520 4680 1580 4690
rect 1520 4660 1530 4680
rect 1570 4660 1580 4680
rect 1520 4650 1580 4660
rect 1740 4680 1800 4690
rect 1740 4660 1750 4680
rect 1790 4660 1800 4680
rect 1740 4650 1800 4660
rect 1910 4680 1970 4690
rect 1910 4660 1920 4680
rect 1960 4660 1970 4680
rect 1910 4650 1970 4660
rect 2080 4680 2140 4690
rect 2080 4660 2090 4680
rect 2130 4660 2140 4680
rect 2080 4650 2140 4660
rect 2250 4680 2310 4690
rect 2250 4660 2260 4680
rect 2300 4660 2310 4680
rect 2250 4650 2310 4660
rect 2420 4680 2480 4690
rect 2420 4660 2430 4680
rect 2470 4660 2480 4680
rect 2420 4650 2480 4660
rect 2590 4680 2650 4690
rect 2590 4660 2600 4680
rect 2640 4660 2650 4680
rect 2590 4650 2650 4660
rect 2760 4680 2820 4690
rect 2760 4660 2770 4680
rect 2810 4660 2820 4680
rect 2760 4650 2820 4660
rect 2930 4680 2990 4690
rect 2930 4660 2940 4680
rect 2980 4660 2990 4680
rect 2930 4650 2990 4660
rect 3100 4680 3160 4690
rect 3100 4660 3110 4680
rect 3150 4660 3160 4680
rect 3100 4650 3160 4660
rect 3270 4680 3330 4690
rect 3270 4660 3280 4680
rect 3320 4660 3330 4680
rect 3270 4650 3330 4660
rect -30 2520 70 2530
rect -30 2500 0 2520
rect 40 2500 70 2520
rect 140 2520 240 2530
rect 140 2500 170 2520
rect 210 2500 240 2520
rect 310 2520 410 2530
rect 310 2500 340 2520
rect 380 2500 410 2520
rect 480 2520 580 2530
rect 480 2500 510 2520
rect 550 2500 580 2520
rect 650 2520 750 2530
rect 650 2500 680 2520
rect 720 2500 750 2520
rect 820 2520 920 2530
rect 820 2500 850 2520
rect 890 2500 920 2520
rect 990 2520 1090 2530
rect 990 2500 1020 2520
rect 1060 2500 1090 2520
rect 1160 2520 1260 2530
rect 1160 2500 1190 2520
rect 1230 2500 1260 2520
rect 1330 2520 1430 2530
rect 1330 2500 1360 2520
rect 1400 2500 1430 2520
rect 1500 2520 1600 2530
rect 1500 2500 1530 2520
rect 1570 2500 1600 2520
rect 1720 2520 1820 2530
rect 1720 2500 1750 2520
rect 1790 2500 1820 2520
rect 1890 2520 1990 2530
rect 1890 2500 1920 2520
rect 1960 2500 1990 2520
rect 2060 2520 2160 2530
rect 2060 2500 2090 2520
rect 2130 2500 2160 2520
rect 2230 2520 2330 2530
rect 2230 2500 2260 2520
rect 2300 2500 2330 2520
rect 2400 2520 2500 2530
rect 2400 2500 2430 2520
rect 2470 2500 2500 2520
rect 2570 2520 2670 2530
rect 2570 2500 2600 2520
rect 2640 2500 2670 2520
rect 2740 2520 2840 2530
rect 2740 2500 2770 2520
rect 2810 2500 2840 2520
rect 2910 2520 3010 2530
rect 2910 2500 2940 2520
rect 2980 2500 3010 2520
rect 3080 2520 3180 2530
rect 3080 2500 3110 2520
rect 3150 2500 3180 2520
rect 3250 2520 3350 2530
rect 3250 2500 3280 2520
rect 3320 2500 3350 2520
<< nsubdiff >>
rect -270 5210 -230 5220
rect -270 5170 -260 5210
rect -240 5170 -230 5210
rect -270 5160 -230 5170
rect 3550 5210 3590 5220
rect 3550 5170 3560 5210
rect 3580 5170 3590 5210
rect 3550 5160 3590 5170
rect 1370 5100 1430 5120
rect 1370 5080 1390 5100
rect 1410 5080 1430 5100
rect 1370 5060 1430 5080
rect 1890 5100 1950 5120
rect 1890 5080 1910 5100
rect 1930 5080 1950 5100
rect 1890 5060 1950 5080
rect -270 5010 -230 5020
rect -270 4970 -260 5010
rect -240 4970 -230 5010
rect -270 4960 -230 4970
rect 3550 5010 3590 5020
rect 3550 4970 3560 5010
rect 3580 4970 3590 5010
rect 3550 4960 3590 4970
<< psubdiffcont >>
rect 0 7660 40 7680
rect 170 7660 210 7680
rect 340 7660 380 7680
rect 510 7660 550 7680
rect 680 7660 720 7680
rect 850 7660 890 7680
rect 1020 7660 1060 7680
rect 1190 7660 1230 7680
rect 1360 7660 1400 7680
rect 1530 7660 1570 7680
rect 1750 7660 1790 7680
rect 1920 7660 1960 7680
rect 2090 7660 2130 7680
rect 2260 7660 2300 7680
rect 2430 7660 2470 7680
rect 2600 7660 2640 7680
rect 2770 7660 2810 7680
rect 2940 7660 2980 7680
rect 3110 7660 3150 7680
rect 3280 7660 3320 7680
rect 0 5500 40 5520
rect 170 5500 210 5520
rect 340 5500 380 5520
rect 510 5500 550 5520
rect 680 5500 720 5520
rect 850 5500 890 5520
rect 1020 5500 1060 5520
rect 1190 5500 1230 5520
rect 1360 5500 1400 5520
rect 1530 5500 1570 5520
rect 1750 5500 1790 5520
rect 1920 5500 1960 5520
rect 2090 5500 2130 5520
rect 2260 5500 2300 5520
rect 2430 5500 2470 5520
rect 2600 5500 2640 5520
rect 2770 5500 2810 5520
rect 2940 5500 2980 5520
rect 3110 5500 3150 5520
rect 3280 5500 3320 5520
rect 0 4660 40 4680
rect 170 4660 210 4680
rect 340 4660 380 4680
rect 510 4660 550 4680
rect 680 4660 720 4680
rect 850 4660 890 4680
rect 1020 4660 1060 4680
rect 1190 4660 1230 4680
rect 1360 4660 1400 4680
rect 1530 4660 1570 4680
rect 1750 4660 1790 4680
rect 1920 4660 1960 4680
rect 2090 4660 2130 4680
rect 2260 4660 2300 4680
rect 2430 4660 2470 4680
rect 2600 4660 2640 4680
rect 2770 4660 2810 4680
rect 2940 4660 2980 4680
rect 3110 4660 3150 4680
rect 3280 4660 3320 4680
rect 0 2500 40 2520
rect 170 2500 210 2520
rect 340 2500 380 2520
rect 510 2500 550 2520
rect 680 2500 720 2520
rect 850 2500 890 2520
rect 1020 2500 1060 2520
rect 1190 2500 1230 2520
rect 1360 2500 1400 2520
rect 1530 2500 1570 2520
rect 1750 2500 1790 2520
rect 1920 2500 1960 2520
rect 2090 2500 2130 2520
rect 2260 2500 2300 2520
rect 2430 2500 2470 2520
rect 2600 2500 2640 2520
rect 2770 2500 2810 2520
rect 2940 2500 2980 2520
rect 3110 2500 3150 2520
rect 3280 2500 3320 2520
<< nsubdiffcont >>
rect -260 5170 -240 5210
rect 3560 5170 3580 5210
rect 1390 5080 1410 5100
rect 1910 5080 1930 5100
rect -260 4970 -240 5010
rect 3560 4970 3580 5010
<< poly >>
rect -90 7660 -50 7670
rect -90 7640 -80 7660
rect -60 7640 -50 7660
rect -90 7630 -50 7640
rect -70 7610 -50 7630
rect 3370 7660 3410 7670
rect 3370 7640 3380 7660
rect 3400 7640 3410 7660
rect 3370 7630 3410 7640
rect 3370 7610 3390 7630
rect -70 7590 -30 7610
rect -340 6660 -300 6670
rect -340 6640 -330 6660
rect -310 6640 -300 6660
rect -340 6630 -300 6640
rect -340 6570 -320 6630
rect -50 6610 -30 7590
rect 70 7120 90 7610
rect 120 7120 140 7610
rect 70 7100 140 7120
rect 70 6610 90 7100
rect 120 6610 140 7100
rect 240 7120 260 7610
rect 290 7120 310 7610
rect 240 7100 310 7120
rect 240 6610 260 7100
rect 290 6610 310 7100
rect 410 7120 430 7610
rect 460 7120 480 7610
rect 410 7100 480 7120
rect 410 6610 430 7100
rect 460 6610 480 7100
rect 580 7120 600 7610
rect 630 7120 650 7610
rect 580 7100 650 7120
rect 580 6610 600 7100
rect 630 6610 650 7100
rect 750 7120 770 7610
rect 800 7120 820 7610
rect 750 7100 820 7120
rect 750 6610 770 7100
rect 800 6610 820 7100
rect 920 7120 940 7610
rect 970 7120 990 7610
rect 920 7100 990 7120
rect 920 6610 940 7100
rect 970 6610 990 7100
rect 1090 7120 1110 7610
rect 1140 7120 1160 7610
rect 1090 7100 1160 7120
rect 1090 6610 1110 7100
rect 1140 6610 1160 7100
rect 1260 7120 1280 7610
rect 1310 7120 1330 7610
rect 1260 7100 1330 7120
rect 1260 6610 1280 7100
rect 1310 6610 1330 7100
rect 1430 7120 1450 7610
rect 1480 7120 1500 7610
rect 1430 7100 1500 7120
rect 1430 6610 1450 7100
rect 1480 6610 1500 7100
rect 1600 7120 1620 7610
rect 1700 7120 1720 7610
rect 1600 7100 1720 7120
rect 1600 6610 1620 7100
rect 1700 6610 1720 7100
rect 1820 7120 1840 7610
rect 1870 7120 1890 7610
rect 1820 7100 1890 7120
rect 1820 6610 1840 7100
rect 1870 6610 1890 7100
rect 1990 7120 2010 7610
rect 2040 7120 2060 7610
rect 1990 7100 2060 7120
rect 1990 6610 2010 7100
rect 2040 6610 2060 7100
rect 2160 7120 2180 7610
rect 2210 7120 2230 7610
rect 2160 7100 2230 7120
rect 2160 6610 2180 7100
rect 2210 6610 2230 7100
rect 2330 7120 2350 7610
rect 2380 7120 2400 7610
rect 2330 7100 2400 7120
rect 2330 6610 2350 7100
rect 2380 6610 2400 7100
rect 2500 7120 2520 7610
rect 2550 7120 2570 7610
rect 2500 7100 2570 7120
rect 2500 6610 2520 7100
rect 2550 6610 2570 7100
rect 2670 7120 2690 7610
rect 2720 7120 2740 7610
rect 2670 7100 2740 7120
rect 2670 6610 2690 7100
rect 2720 6610 2740 7100
rect 2840 7120 2860 7610
rect 2890 7120 2910 7610
rect 2840 7100 2910 7120
rect 2840 6610 2860 7100
rect 2890 6610 2910 7100
rect 3010 7120 3030 7610
rect 3060 7120 3080 7610
rect 3010 7100 3080 7120
rect 3010 6610 3030 7100
rect 3060 6610 3080 7100
rect 3180 7120 3200 7610
rect 3230 7120 3250 7610
rect 3180 7100 3250 7120
rect 3180 6610 3200 7100
rect 3230 6610 3250 7100
rect 3350 7590 3390 7610
rect 3350 6610 3370 7590
rect 3620 6660 3660 6670
rect 3620 6640 3630 6660
rect 3650 6640 3660 6660
rect 3620 6630 3660 6640
rect 3640 6570 3660 6630
rect -340 6550 -310 6570
rect -330 6070 -310 6550
rect -110 6070 -90 6570
rect -330 5530 -310 6030
rect -110 5550 -90 6030
rect -50 5570 -30 6570
rect 70 6080 90 6570
rect 120 6080 140 6570
rect 70 6060 140 6080
rect 70 5570 90 6060
rect 120 5570 140 6060
rect 240 6080 260 6570
rect 290 6080 310 6570
rect 240 6060 310 6080
rect 240 5570 260 6060
rect 290 5570 310 6060
rect 410 6080 430 6570
rect 460 6080 480 6570
rect 410 6060 480 6080
rect 410 5570 430 6060
rect 460 5570 480 6060
rect 580 6080 600 6570
rect 630 6080 650 6570
rect 580 6060 650 6080
rect 580 5570 600 6060
rect 630 5570 650 6060
rect 750 6080 770 6570
rect 800 6080 820 6570
rect 750 6060 820 6080
rect 750 5570 770 6060
rect 800 5570 820 6060
rect 920 6080 940 6570
rect 970 6080 990 6570
rect 920 6060 990 6080
rect 920 5570 940 6060
rect 970 5570 990 6060
rect 1090 6080 1110 6570
rect 1140 6080 1160 6570
rect 1090 6060 1160 6080
rect 1090 5570 1110 6060
rect 1140 5570 1160 6060
rect 1260 6080 1280 6570
rect 1310 6080 1330 6570
rect 1260 6060 1330 6080
rect 1260 5570 1280 6060
rect 1310 5570 1330 6060
rect 1430 6080 1450 6570
rect 1480 6080 1500 6570
rect 1430 6060 1500 6080
rect 1430 5570 1450 6060
rect 1480 5570 1500 6060
rect 1600 6080 1620 6570
rect 1700 6080 1720 6570
rect 1600 6060 1720 6080
rect 1600 5570 1620 6060
rect -110 5530 -80 5550
rect -100 5470 -80 5530
rect -120 5460 -80 5470
rect -120 5440 -110 5460
rect -90 5440 -80 5460
rect -120 5430 -80 5440
rect -50 5360 -30 5460
rect 70 5420 90 5460
rect 120 5420 140 5460
rect 70 5400 140 5420
rect 70 5360 90 5400
rect 120 5360 140 5400
rect 240 5420 260 5460
rect 290 5420 310 5460
rect 240 5400 310 5420
rect 240 5360 260 5400
rect 290 5360 310 5400
rect 410 5420 430 5460
rect 460 5420 480 5460
rect 410 5400 480 5420
rect 410 5360 430 5400
rect 460 5360 480 5400
rect 580 5420 600 5460
rect 630 5420 650 5460
rect 580 5400 650 5420
rect 580 5360 600 5400
rect 630 5360 650 5400
rect 750 5420 770 5460
rect 800 5420 820 5460
rect 750 5400 820 5420
rect 750 5360 770 5400
rect 800 5360 820 5400
rect 920 5420 940 5460
rect 970 5420 990 5460
rect 920 5400 990 5420
rect 920 5360 940 5400
rect 970 5360 990 5400
rect 1090 5420 1110 5460
rect 1140 5420 1160 5460
rect 1090 5400 1160 5420
rect 1090 5360 1110 5400
rect 1140 5360 1160 5400
rect 1260 5420 1280 5460
rect 1310 5420 1330 5460
rect 1260 5400 1330 5420
rect 1260 5360 1280 5400
rect 1310 5360 1330 5400
rect 1430 5420 1450 5460
rect 1480 5420 1500 5460
rect 1430 5400 1500 5420
rect 1430 5360 1450 5400
rect 1480 5360 1500 5400
rect 1600 5420 1620 5460
rect 1650 5420 1670 6060
rect 1700 5570 1720 6060
rect 1820 6080 1840 6570
rect 1870 6080 1890 6570
rect 1820 6060 1890 6080
rect 1820 5570 1840 6060
rect 1870 5570 1890 6060
rect 1990 6080 2010 6570
rect 2040 6080 2060 6570
rect 1990 6060 2060 6080
rect 1990 5570 2010 6060
rect 2040 5570 2060 6060
rect 2160 6080 2180 6570
rect 2210 6080 2230 6570
rect 2160 6060 2230 6080
rect 2160 5570 2180 6060
rect 2210 5570 2230 6060
rect 2330 6080 2350 6570
rect 2380 6080 2400 6570
rect 2330 6060 2400 6080
rect 2330 5570 2350 6060
rect 2380 5570 2400 6060
rect 2500 6080 2520 6570
rect 2550 6080 2570 6570
rect 2500 6060 2570 6080
rect 2500 5570 2520 6060
rect 2550 5570 2570 6060
rect 2670 6080 2690 6570
rect 2720 6080 2740 6570
rect 2670 6060 2740 6080
rect 2670 5570 2690 6060
rect 2720 5570 2740 6060
rect 2840 6080 2860 6570
rect 2890 6080 2910 6570
rect 2840 6060 2910 6080
rect 2840 5570 2860 6060
rect 2890 5570 2910 6060
rect 3010 6080 3030 6570
rect 3060 6080 3080 6570
rect 3010 6060 3080 6080
rect 3010 5570 3030 6060
rect 3060 5570 3080 6060
rect 3180 6080 3200 6570
rect 3230 6080 3250 6570
rect 3180 6060 3250 6080
rect 3180 5570 3200 6060
rect 3230 5570 3250 6060
rect 3350 5570 3370 6570
rect 3410 6070 3430 6570
rect 3630 6550 3660 6570
rect 3630 6070 3650 6550
rect 3410 5550 3430 6030
rect 3400 5530 3430 5550
rect 3630 5530 3650 6030
rect 3400 5470 3420 5530
rect 3400 5460 3440 5470
rect 1700 5420 1720 5460
rect 1600 5400 1720 5420
rect 1600 5360 1630 5400
rect 1610 5300 1630 5360
rect -230 5290 -190 5300
rect -230 5270 -220 5290
rect -200 5280 -190 5290
rect 50 5290 90 5300
rect 50 5280 60 5290
rect -200 5270 -170 5280
rect -230 5260 -170 5270
rect 30 5270 60 5280
rect 80 5280 90 5290
rect 330 5290 370 5300
rect 330 5280 340 5290
rect 80 5270 110 5280
rect 30 5260 110 5270
rect 310 5270 340 5280
rect 360 5280 370 5290
rect 610 5290 650 5300
rect 610 5280 620 5290
rect 360 5270 390 5280
rect 310 5260 390 5270
rect 590 5270 620 5280
rect 640 5280 650 5290
rect 890 5290 930 5300
rect 890 5280 900 5290
rect 640 5270 670 5280
rect 590 5260 670 5270
rect 870 5270 900 5280
rect 920 5280 930 5290
rect 1170 5290 1210 5300
rect 1170 5280 1180 5290
rect 920 5270 950 5280
rect 870 5260 950 5270
rect 1150 5270 1180 5280
rect 1200 5280 1210 5290
rect 1580 5290 1630 5300
rect 1200 5270 1230 5280
rect 1150 5260 1230 5270
rect 1580 5270 1590 5290
rect 1610 5270 1630 5290
rect 1580 5260 1630 5270
rect 1690 5360 1720 5400
rect 1820 5420 1840 5460
rect 1870 5420 1890 5460
rect 1820 5400 1890 5420
rect 1820 5360 1840 5400
rect 1870 5360 1890 5400
rect 1990 5420 2010 5460
rect 2040 5420 2060 5460
rect 1990 5400 2060 5420
rect 1990 5360 2010 5400
rect 2040 5360 2060 5400
rect 2160 5420 2180 5460
rect 2210 5420 2230 5460
rect 2160 5400 2230 5420
rect 2160 5360 2180 5400
rect 2210 5360 2230 5400
rect 2330 5420 2350 5460
rect 2380 5420 2400 5460
rect 2330 5400 2400 5420
rect 2330 5360 2350 5400
rect 2380 5360 2400 5400
rect 2500 5420 2520 5460
rect 2550 5420 2570 5460
rect 2500 5400 2570 5420
rect 2500 5360 2520 5400
rect 2550 5360 2570 5400
rect 2670 5420 2690 5460
rect 2720 5420 2740 5460
rect 2670 5400 2740 5420
rect 2670 5360 2690 5400
rect 2720 5360 2740 5400
rect 2840 5420 2860 5460
rect 2890 5420 2910 5460
rect 2840 5400 2910 5420
rect 2840 5360 2860 5400
rect 2890 5360 2910 5400
rect 3010 5420 3030 5460
rect 3060 5420 3080 5460
rect 3010 5400 3080 5420
rect 3010 5360 3030 5400
rect 3060 5360 3080 5400
rect 3180 5420 3200 5460
rect 3230 5420 3250 5460
rect 3180 5400 3250 5420
rect 3180 5360 3200 5400
rect 3230 5360 3250 5400
rect 3350 5360 3370 5460
rect 3400 5440 3410 5460
rect 3430 5440 3440 5460
rect 3400 5430 3440 5440
rect 1690 5300 1710 5360
rect 1690 5290 1740 5300
rect 1690 5270 1710 5290
rect 1730 5270 1740 5290
rect 2110 5290 2150 5300
rect 2110 5280 2120 5290
rect 1690 5260 1740 5270
rect 2090 5270 2120 5280
rect 2140 5280 2150 5290
rect 2390 5290 2430 5300
rect 2390 5280 2400 5290
rect 2140 5270 2170 5280
rect 2090 5260 2170 5270
rect 2370 5270 2400 5280
rect 2420 5280 2430 5290
rect 2670 5290 2710 5300
rect 2670 5280 2680 5290
rect 2420 5270 2450 5280
rect 2370 5260 2450 5270
rect 2650 5270 2680 5280
rect 2700 5280 2710 5290
rect 2950 5290 2990 5300
rect 2950 5280 2960 5290
rect 2700 5270 2730 5280
rect 2650 5260 2730 5270
rect 2930 5270 2960 5280
rect 2980 5280 2990 5290
rect 3230 5290 3270 5300
rect 3230 5280 3240 5290
rect 2980 5270 3010 5280
rect 2930 5260 3010 5270
rect 3210 5270 3240 5280
rect 3260 5280 3270 5290
rect 3510 5290 3550 5300
rect 3510 5280 3520 5290
rect 3260 5270 3290 5280
rect 3210 5260 3290 5270
rect 3490 5270 3520 5280
rect 3540 5270 3550 5290
rect 3490 5260 3550 5270
rect -190 5240 -90 5260
rect -50 5240 50 5260
rect 90 5240 190 5260
rect 230 5240 330 5260
rect 370 5240 470 5260
rect 510 5240 610 5260
rect 650 5240 750 5260
rect 790 5240 890 5260
rect 930 5240 1030 5260
rect 1070 5240 1170 5260
rect 1210 5240 1310 5260
rect 2010 5240 2110 5260
rect 2150 5240 2250 5260
rect 2290 5240 2390 5260
rect 2430 5240 2530 5260
rect 2570 5240 2670 5260
rect 2710 5240 2810 5260
rect 2850 5240 2950 5260
rect 2990 5240 3090 5260
rect 3130 5240 3230 5260
rect 3270 5240 3370 5260
rect 3410 5240 3510 5260
rect -190 5120 -90 5140
rect -50 5120 50 5140
rect 90 5120 190 5140
rect 230 5120 330 5140
rect 370 5120 470 5140
rect 510 5120 610 5140
rect 650 5120 750 5140
rect 790 5120 890 5140
rect 930 5120 1030 5140
rect 1070 5120 1170 5140
rect -190 5040 -90 5060
rect -50 5040 50 5060
rect 90 5040 190 5060
rect 230 5040 330 5060
rect 370 5040 470 5060
rect 510 5040 610 5060
rect 650 5040 750 5060
rect 790 5040 890 5060
rect 930 5040 1030 5060
rect 1070 5040 1170 5060
rect 1210 5120 1310 5140
rect 1210 5040 1310 5060
rect 2010 5120 2110 5140
rect 2010 5040 2110 5060
rect 2150 5120 2250 5140
rect 2290 5120 2390 5140
rect 2430 5120 2530 5140
rect 2570 5120 2670 5140
rect 2710 5120 2810 5140
rect 2850 5120 2950 5140
rect 2990 5120 3090 5140
rect 3130 5120 3230 5140
rect 3270 5120 3370 5140
rect 3410 5120 3510 5140
rect 2150 5040 2250 5060
rect 2290 5040 2390 5060
rect 2430 5040 2530 5060
rect 2570 5040 2670 5060
rect 2710 5040 2810 5060
rect 2850 5040 2950 5060
rect 2990 5040 3090 5060
rect 3130 5040 3230 5060
rect 3270 5040 3370 5060
rect 3410 5040 3510 5060
rect -190 4920 -90 4940
rect -50 4920 50 4940
rect 90 4920 190 4940
rect 230 4920 330 4940
rect 370 4920 470 4940
rect 510 4920 610 4940
rect 650 4920 750 4940
rect 790 4920 890 4940
rect 930 4920 1030 4940
rect 1070 4920 1170 4940
rect 1210 4920 1310 4940
rect 2010 4920 2110 4940
rect 2150 4920 2250 4940
rect 2290 4920 2390 4940
rect 2430 4920 2530 4940
rect 2570 4920 2670 4940
rect 2710 4920 2810 4940
rect 2850 4920 2950 4940
rect 2990 4920 3090 4940
rect 3130 4920 3230 4940
rect 3270 4920 3370 4940
rect 3410 4920 3510 4940
rect -230 4910 -170 4920
rect -230 4890 -220 4910
rect -200 4900 -170 4910
rect 30 4910 110 4920
rect 30 4900 60 4910
rect -200 4890 -190 4900
rect -230 4880 -190 4890
rect 50 4890 60 4900
rect 80 4900 110 4910
rect 310 4910 390 4920
rect 310 4900 340 4910
rect 80 4890 90 4900
rect 50 4880 90 4890
rect 330 4890 340 4900
rect 360 4900 390 4910
rect 590 4910 670 4920
rect 590 4900 620 4910
rect 360 4890 370 4900
rect 330 4880 370 4890
rect 610 4890 620 4900
rect 640 4900 670 4910
rect 870 4910 950 4920
rect 870 4900 900 4910
rect 640 4890 650 4900
rect 610 4880 650 4890
rect 890 4890 900 4900
rect 920 4900 950 4910
rect 1150 4910 1230 4920
rect 1150 4900 1180 4910
rect 920 4890 930 4900
rect 890 4880 930 4890
rect 1170 4890 1180 4900
rect 1200 4900 1230 4910
rect 1580 4910 1630 4920
rect 1200 4890 1210 4900
rect 1170 4880 1210 4890
rect 1580 4890 1590 4910
rect 1610 4890 1630 4910
rect 1580 4880 1630 4890
rect 1610 4820 1630 4880
rect -120 4740 -80 4750
rect -120 4720 -110 4740
rect -90 4720 -80 4740
rect -50 4720 -30 4820
rect 70 4780 90 4820
rect 120 4780 140 4820
rect 70 4760 140 4780
rect 70 4720 90 4760
rect 120 4720 140 4760
rect 240 4780 260 4820
rect 290 4780 310 4820
rect 240 4760 310 4780
rect 240 4720 260 4760
rect 290 4720 310 4760
rect 410 4780 430 4820
rect 460 4780 480 4820
rect 410 4760 480 4780
rect 410 4720 430 4760
rect 460 4720 480 4760
rect 580 4780 600 4820
rect 630 4780 650 4820
rect 580 4760 650 4780
rect 580 4720 600 4760
rect 630 4720 650 4760
rect 750 4780 770 4820
rect 800 4780 820 4820
rect 750 4760 820 4780
rect 750 4720 770 4760
rect 800 4720 820 4760
rect 920 4780 940 4820
rect 970 4780 990 4820
rect 920 4760 990 4780
rect 920 4720 940 4760
rect 970 4720 990 4760
rect 1090 4780 1110 4820
rect 1140 4780 1160 4820
rect 1090 4760 1160 4780
rect 1090 4720 1110 4760
rect 1140 4720 1160 4760
rect 1260 4780 1280 4820
rect 1310 4780 1330 4820
rect 1260 4760 1330 4780
rect 1260 4720 1280 4760
rect 1310 4720 1330 4760
rect 1430 4780 1450 4820
rect 1480 4780 1500 4820
rect 1430 4760 1500 4780
rect 1430 4720 1450 4760
rect 1480 4720 1500 4760
rect 1600 4780 1630 4820
rect 1690 4910 1740 4920
rect 1690 4890 1710 4910
rect 1730 4890 1740 4910
rect 2090 4910 2170 4920
rect 2090 4900 2120 4910
rect 1690 4880 1740 4890
rect 2110 4890 2120 4900
rect 2140 4900 2170 4910
rect 2370 4910 2450 4920
rect 2370 4900 2400 4910
rect 2140 4890 2150 4900
rect 2110 4880 2150 4890
rect 2390 4890 2400 4900
rect 2420 4900 2450 4910
rect 2650 4910 2730 4920
rect 2650 4900 2680 4910
rect 2420 4890 2430 4900
rect 2390 4880 2430 4890
rect 2670 4890 2680 4900
rect 2700 4900 2730 4910
rect 2930 4910 3010 4920
rect 2930 4900 2960 4910
rect 2700 4890 2710 4900
rect 2670 4880 2710 4890
rect 2950 4890 2960 4900
rect 2980 4900 3010 4910
rect 3210 4910 3290 4920
rect 3210 4900 3240 4910
rect 2980 4890 2990 4900
rect 2950 4880 2990 4890
rect 3230 4890 3240 4900
rect 3260 4900 3290 4910
rect 3490 4910 3550 4920
rect 3490 4900 3520 4910
rect 3260 4890 3270 4900
rect 3230 4880 3270 4890
rect 3510 4890 3520 4900
rect 3540 4890 3550 4910
rect 3510 4880 3550 4890
rect 1690 4820 1710 4880
rect 1690 4780 1720 4820
rect 1600 4760 1720 4780
rect 1600 4720 1620 4760
rect -120 4710 -80 4720
rect -100 4650 -80 4710
rect -330 4150 -310 4650
rect -110 4630 -80 4650
rect -110 4150 -90 4630
rect -330 3630 -310 4110
rect -340 3610 -310 3630
rect -110 3610 -90 4110
rect -50 3610 -30 4610
rect 70 4120 90 4610
rect 120 4120 140 4610
rect 70 4100 140 4120
rect 70 3610 90 4100
rect 120 3610 140 4100
rect 240 4120 260 4610
rect 290 4120 310 4610
rect 240 4100 310 4120
rect 240 3610 260 4100
rect 290 3610 310 4100
rect 410 4120 430 4610
rect 460 4120 480 4610
rect 410 4100 480 4120
rect 410 3610 430 4100
rect 460 3610 480 4100
rect 580 4120 600 4610
rect 630 4120 650 4610
rect 580 4100 650 4120
rect 580 3610 600 4100
rect 630 3610 650 4100
rect 750 4120 770 4610
rect 800 4120 820 4610
rect 750 4100 820 4120
rect 750 3610 770 4100
rect 800 3610 820 4100
rect 920 4120 940 4610
rect 970 4120 990 4610
rect 920 4100 990 4120
rect 920 3610 940 4100
rect 970 3610 990 4100
rect 1090 4120 1110 4610
rect 1140 4120 1160 4610
rect 1090 4100 1160 4120
rect 1090 3610 1110 4100
rect 1140 3610 1160 4100
rect 1260 4120 1280 4610
rect 1310 4120 1330 4610
rect 1260 4100 1330 4120
rect 1260 3610 1280 4100
rect 1310 3610 1330 4100
rect 1430 4120 1450 4610
rect 1480 4120 1500 4610
rect 1430 4100 1500 4120
rect 1430 3610 1450 4100
rect 1480 3610 1500 4100
rect 1600 4120 1620 4610
rect 1650 4120 1670 4760
rect 1700 4720 1720 4760
rect 1820 4780 1840 4820
rect 1870 4780 1890 4820
rect 1820 4760 1890 4780
rect 1820 4720 1840 4760
rect 1870 4720 1890 4760
rect 1990 4780 2010 4820
rect 2040 4780 2060 4820
rect 1990 4760 2060 4780
rect 1990 4720 2010 4760
rect 2040 4720 2060 4760
rect 2160 4780 2180 4820
rect 2210 4780 2230 4820
rect 2160 4760 2230 4780
rect 2160 4720 2180 4760
rect 2210 4720 2230 4760
rect 2330 4780 2350 4820
rect 2380 4780 2400 4820
rect 2330 4760 2400 4780
rect 2330 4720 2350 4760
rect 2380 4720 2400 4760
rect 2500 4780 2520 4820
rect 2550 4780 2570 4820
rect 2500 4760 2570 4780
rect 2500 4720 2520 4760
rect 2550 4720 2570 4760
rect 2670 4780 2690 4820
rect 2720 4780 2740 4820
rect 2670 4760 2740 4780
rect 2670 4720 2690 4760
rect 2720 4720 2740 4760
rect 2840 4780 2860 4820
rect 2890 4780 2910 4820
rect 2840 4760 2910 4780
rect 2840 4720 2860 4760
rect 2890 4720 2910 4760
rect 3010 4780 3030 4820
rect 3060 4780 3080 4820
rect 3010 4760 3080 4780
rect 3010 4720 3030 4760
rect 3060 4720 3080 4760
rect 3180 4780 3200 4820
rect 3230 4780 3250 4820
rect 3180 4760 3250 4780
rect 3180 4720 3200 4760
rect 3230 4720 3250 4760
rect 3350 4720 3370 4820
rect 3400 4740 3440 4750
rect 3400 4720 3410 4740
rect 3430 4720 3440 4740
rect 3400 4710 3440 4720
rect 3400 4650 3420 4710
rect 3400 4630 3430 4650
rect 1700 4120 1720 4610
rect 1600 4100 1720 4120
rect 1600 3610 1620 4100
rect 1700 3610 1720 4100
rect 1820 4120 1840 4610
rect 1870 4120 1890 4610
rect 1820 4100 1890 4120
rect 1820 3610 1840 4100
rect 1870 3610 1890 4100
rect 1990 4120 2010 4610
rect 2040 4120 2060 4610
rect 1990 4100 2060 4120
rect 1990 3610 2010 4100
rect 2040 3610 2060 4100
rect 2160 4120 2180 4610
rect 2210 4120 2230 4610
rect 2160 4100 2230 4120
rect 2160 3610 2180 4100
rect 2210 3610 2230 4100
rect 2330 4120 2350 4610
rect 2380 4120 2400 4610
rect 2330 4100 2400 4120
rect 2330 3610 2350 4100
rect 2380 3610 2400 4100
rect 2500 4120 2520 4610
rect 2550 4120 2570 4610
rect 2500 4100 2570 4120
rect 2500 3610 2520 4100
rect 2550 3610 2570 4100
rect 2670 4120 2690 4610
rect 2720 4120 2740 4610
rect 2670 4100 2740 4120
rect 2670 3610 2690 4100
rect 2720 3610 2740 4100
rect 2840 4120 2860 4610
rect 2890 4120 2910 4610
rect 2840 4100 2910 4120
rect 2840 3610 2860 4100
rect 2890 3610 2910 4100
rect 3010 4120 3030 4610
rect 3060 4120 3080 4610
rect 3010 4100 3080 4120
rect 3010 3610 3030 4100
rect 3060 3610 3080 4100
rect 3180 4120 3200 4610
rect 3230 4120 3250 4610
rect 3180 4100 3250 4120
rect 3180 3610 3200 4100
rect 3230 3610 3250 4100
rect 3350 3610 3370 4610
rect 3410 4150 3430 4630
rect 3630 4150 3650 4650
rect 3410 3610 3430 4110
rect 3630 3630 3650 4110
rect 3630 3610 3660 3630
rect -340 3550 -320 3610
rect -340 3540 -300 3550
rect -340 3520 -330 3540
rect -310 3520 -300 3540
rect -340 3510 -300 3520
rect -50 2590 -30 3570
rect -70 2570 -30 2590
rect 70 3080 90 3570
rect 120 3080 140 3570
rect 70 3060 140 3080
rect 70 2570 90 3060
rect 120 2570 140 3060
rect 240 3080 260 3570
rect 290 3080 310 3570
rect 240 3060 310 3080
rect 240 2570 260 3060
rect 290 2570 310 3060
rect 410 3080 430 3570
rect 460 3080 480 3570
rect 410 3060 480 3080
rect 410 2570 430 3060
rect 460 2570 480 3060
rect 580 3080 600 3570
rect 630 3080 650 3570
rect 580 3060 650 3080
rect 580 2570 600 3060
rect 630 2570 650 3060
rect 750 3080 770 3570
rect 800 3080 820 3570
rect 750 3060 820 3080
rect 750 2570 770 3060
rect 800 2570 820 3060
rect 920 3080 940 3570
rect 970 3080 990 3570
rect 920 3060 990 3080
rect 920 2570 940 3060
rect 970 2570 990 3060
rect 1090 3080 1110 3570
rect 1140 3080 1160 3570
rect 1090 3060 1160 3080
rect 1090 2570 1110 3060
rect 1140 2570 1160 3060
rect 1260 3080 1280 3570
rect 1310 3080 1330 3570
rect 1260 3060 1330 3080
rect 1260 2570 1280 3060
rect 1310 2570 1330 3060
rect 1430 3080 1450 3570
rect 1480 3080 1500 3570
rect 1430 3060 1500 3080
rect 1430 2570 1450 3060
rect 1480 2570 1500 3060
rect 1600 3080 1620 3570
rect 1700 3080 1720 3570
rect 1600 3060 1720 3080
rect 1600 2570 1620 3060
rect 1700 2570 1720 3060
rect 1820 3080 1840 3570
rect 1870 3080 1890 3570
rect 1820 3060 1890 3080
rect 1820 2570 1840 3060
rect 1870 2570 1890 3060
rect 1990 3080 2010 3570
rect 2040 3080 2060 3570
rect 1990 3060 2060 3080
rect 1990 2570 2010 3060
rect 2040 2570 2060 3060
rect 2160 3080 2180 3570
rect 2210 3080 2230 3570
rect 2160 3060 2230 3080
rect 2160 2570 2180 3060
rect 2210 2570 2230 3060
rect 2330 3080 2350 3570
rect 2380 3080 2400 3570
rect 2330 3060 2400 3080
rect 2330 2570 2350 3060
rect 2380 2570 2400 3060
rect 2500 3080 2520 3570
rect 2550 3080 2570 3570
rect 2500 3060 2570 3080
rect 2500 2570 2520 3060
rect 2550 2570 2570 3060
rect 2670 3080 2690 3570
rect 2720 3080 2740 3570
rect 2670 3060 2740 3080
rect 2670 2570 2690 3060
rect 2720 2570 2740 3060
rect 2840 3080 2860 3570
rect 2890 3080 2910 3570
rect 2840 3060 2910 3080
rect 2840 2570 2860 3060
rect 2890 2570 2910 3060
rect 3010 3080 3030 3570
rect 3060 3080 3080 3570
rect 3010 3060 3080 3080
rect 3010 2570 3030 3060
rect 3060 2570 3080 3060
rect 3180 3080 3200 3570
rect 3230 3080 3250 3570
rect 3180 3060 3250 3080
rect 3180 2570 3200 3060
rect 3230 2570 3250 3060
rect 3350 2590 3370 3570
rect 3640 3550 3660 3610
rect 3620 3540 3660 3550
rect 3620 3520 3630 3540
rect 3650 3520 3660 3540
rect 3620 3510 3660 3520
rect 3350 2570 3390 2590
rect -70 2550 -50 2570
rect -90 2540 -50 2550
rect -90 2520 -80 2540
rect -60 2520 -50 2540
rect -90 2510 -50 2520
rect 3370 2550 3390 2570
rect 3370 2540 3410 2550
rect 3370 2520 3380 2540
rect 3400 2520 3410 2540
rect 3370 2510 3410 2520
<< polycont >>
rect -80 7640 -60 7660
rect 3380 7640 3400 7660
rect -330 6640 -310 6660
rect 3630 6640 3650 6660
rect -110 5440 -90 5460
rect -220 5270 -200 5290
rect 60 5270 80 5290
rect 340 5270 360 5290
rect 620 5270 640 5290
rect 900 5270 920 5290
rect 1180 5270 1200 5290
rect 1590 5270 1610 5290
rect 3410 5440 3430 5460
rect 1710 5270 1730 5290
rect 2120 5270 2140 5290
rect 2400 5270 2420 5290
rect 2680 5270 2700 5290
rect 2960 5270 2980 5290
rect 3240 5270 3260 5290
rect 3520 5270 3540 5290
rect -220 4890 -200 4910
rect 60 4890 80 4910
rect 340 4890 360 4910
rect 620 4890 640 4910
rect 900 4890 920 4910
rect 1180 4890 1200 4910
rect 1590 4890 1610 4910
rect -110 4720 -90 4740
rect 1710 4890 1730 4910
rect 2120 4890 2140 4910
rect 2400 4890 2420 4910
rect 2680 4890 2700 4910
rect 2960 4890 2980 4910
rect 3240 4890 3260 4910
rect 3520 4890 3540 4910
rect 3410 4720 3430 4740
rect -330 3520 -310 3540
rect 3630 3520 3650 3540
rect -80 2520 -60 2540
rect 3380 2520 3400 2540
<< locali >>
rect -90 7660 -50 7670
rect -10 7660 0 7680
rect 40 7660 50 7680
rect 160 7660 170 7680
rect 210 7660 220 7680
rect 330 7660 340 7680
rect 380 7660 390 7680
rect 500 7660 510 7680
rect 550 7660 560 7680
rect 670 7660 680 7680
rect 720 7660 730 7680
rect 840 7660 850 7680
rect 890 7660 900 7680
rect 1010 7660 1020 7680
rect 1060 7660 1070 7680
rect 1180 7660 1190 7680
rect 1230 7660 1240 7680
rect 1350 7660 1360 7680
rect 1400 7660 1410 7680
rect 1520 7660 1530 7680
rect 1570 7660 1580 7680
rect 1740 7660 1750 7680
rect 1790 7660 1800 7680
rect 1910 7660 1920 7680
rect 1960 7660 1970 7680
rect 2080 7660 2090 7680
rect 2130 7660 2140 7680
rect 2250 7660 2260 7680
rect 2300 7660 2310 7680
rect 2420 7660 2430 7680
rect 2470 7660 2480 7680
rect 2590 7660 2600 7680
rect 2640 7660 2650 7680
rect 2760 7660 2770 7680
rect 2810 7660 2820 7680
rect 2930 7660 2940 7680
rect 2980 7660 2990 7680
rect 3100 7660 3110 7680
rect 3150 7660 3160 7680
rect 3270 7660 3280 7680
rect 3320 7660 3330 7680
rect 3370 7660 3410 7670
rect -90 7640 -80 7660
rect -60 7640 3380 7660
rect 3400 7640 3410 7660
rect -90 7630 -50 7640
rect -10 7620 0 7640
rect 40 7620 50 7640
rect -10 7610 50 7620
rect 160 7620 170 7640
rect 210 7620 220 7640
rect 160 7610 220 7620
rect 330 7620 340 7640
rect 380 7620 390 7640
rect 330 7610 390 7620
rect 500 7620 510 7640
rect 550 7620 560 7640
rect 500 7610 560 7620
rect 670 7620 680 7640
rect 720 7620 730 7640
rect 670 7610 730 7620
rect 840 7620 850 7640
rect 890 7620 900 7640
rect 840 7610 900 7620
rect 1010 7620 1020 7640
rect 1060 7620 1070 7640
rect 1010 7610 1070 7620
rect 1180 7620 1190 7640
rect 1230 7620 1240 7640
rect 1180 7610 1240 7620
rect 1350 7620 1360 7640
rect 1400 7620 1410 7640
rect 1350 7610 1410 7620
rect 1520 7620 1530 7640
rect 1570 7620 1580 7640
rect 1520 7610 1580 7620
rect -340 6660 -300 6670
rect -340 6640 -330 6660
rect -310 6640 -200 6660
rect -340 6630 -300 6640
rect -220 6610 -200 6640
rect -240 6600 -180 6610
rect -10 6600 50 6610
rect -240 6580 -230 6600
rect -190 6580 0 6600
rect 40 6580 50 6600
rect -240 6570 -180 6580
rect -10 6570 50 6580
rect 160 6600 220 6610
rect 160 6580 170 6600
rect 210 6580 220 6600
rect 160 6570 220 6580
rect 330 6600 390 6610
rect 330 6580 340 6600
rect 380 6580 390 6600
rect 330 6570 390 6580
rect 500 6600 560 6610
rect 500 6580 510 6600
rect 550 6580 560 6600
rect 500 6570 560 6580
rect 670 6600 730 6610
rect 670 6580 680 6600
rect 720 6580 730 6600
rect 670 6570 730 6580
rect 840 6600 900 6610
rect 840 6580 850 6600
rect 890 6580 900 6600
rect 840 6570 900 6580
rect 1010 6600 1070 6610
rect 1010 6580 1020 6600
rect 1060 6580 1070 6600
rect 1010 6570 1070 6580
rect 1180 6600 1240 6610
rect 1180 6580 1190 6600
rect 1230 6580 1240 6600
rect 1180 6570 1240 6580
rect 1350 6600 1410 6610
rect 1350 6580 1360 6600
rect 1400 6580 1410 6600
rect 1350 6570 1410 6580
rect 1520 6600 1580 6610
rect 1520 6580 1530 6600
rect 1570 6580 1580 6600
rect 1520 6570 1580 6580
rect -240 6060 -180 6070
rect -240 6040 -230 6060
rect -190 6040 -140 6060
rect -240 6030 -180 6040
rect -240 5520 -180 5530
rect -240 5500 -230 5520
rect -190 5500 -180 5520
rect -240 5490 -180 5500
rect -220 5300 -200 5490
rect -160 5310 -140 6040
rect -10 5560 50 5570
rect -10 5540 0 5560
rect 40 5540 50 5560
rect 160 5560 220 5570
rect 160 5540 170 5560
rect 210 5540 220 5560
rect 330 5560 390 5570
rect 330 5540 340 5560
rect 380 5540 390 5560
rect 500 5560 560 5570
rect 500 5540 510 5560
rect 550 5540 560 5560
rect 670 5560 730 5570
rect 670 5540 680 5560
rect 720 5540 730 5560
rect 840 5560 900 5570
rect 840 5540 850 5560
rect 890 5540 900 5560
rect 1010 5560 1070 5570
rect 1010 5540 1020 5560
rect 1060 5540 1070 5560
rect 1180 5560 1240 5570
rect 1180 5540 1190 5560
rect 1230 5540 1240 5560
rect 1350 5560 1410 5570
rect 1350 5540 1360 5560
rect 1400 5540 1410 5560
rect 1520 5560 1580 5570
rect 1520 5540 1530 5560
rect 1570 5540 1580 5560
rect 1650 5540 1670 7640
rect 1740 7620 1750 7640
rect 1790 7620 1800 7640
rect 1740 7610 1800 7620
rect 1910 7620 1920 7640
rect 1960 7620 1970 7640
rect 1910 7610 1970 7620
rect 2080 7620 2090 7640
rect 2130 7620 2140 7640
rect 2080 7610 2140 7620
rect 2250 7620 2260 7640
rect 2300 7620 2310 7640
rect 2250 7610 2310 7620
rect 2420 7620 2430 7640
rect 2470 7620 2480 7640
rect 2420 7610 2480 7620
rect 2590 7620 2600 7640
rect 2640 7620 2650 7640
rect 2590 7610 2650 7620
rect 2760 7620 2770 7640
rect 2810 7620 2820 7640
rect 2760 7610 2820 7620
rect 2930 7620 2940 7640
rect 2980 7620 2990 7640
rect 2930 7610 2990 7620
rect 3100 7620 3110 7640
rect 3150 7620 3160 7640
rect 3100 7610 3160 7620
rect 3270 7620 3280 7640
rect 3320 7620 3330 7640
rect 3370 7630 3410 7640
rect 3270 7610 3330 7620
rect 3620 6660 3660 6670
rect 3520 6640 3630 6660
rect 3650 6640 3660 6660
rect 3520 6610 3540 6640
rect 3620 6630 3660 6640
rect 1740 6600 1800 6610
rect 1740 6580 1750 6600
rect 1790 6580 1800 6600
rect 1740 6570 1800 6580
rect 1910 6600 1970 6610
rect 1910 6580 1920 6600
rect 1960 6580 1970 6600
rect 1910 6570 1970 6580
rect 2080 6600 2140 6610
rect 2080 6580 2090 6600
rect 2130 6580 2140 6600
rect 2080 6570 2140 6580
rect 2250 6600 2310 6610
rect 2250 6580 2260 6600
rect 2300 6580 2310 6600
rect 2250 6570 2310 6580
rect 2420 6600 2480 6610
rect 2420 6580 2430 6600
rect 2470 6580 2480 6600
rect 2420 6570 2480 6580
rect 2590 6600 2650 6610
rect 2590 6580 2600 6600
rect 2640 6580 2650 6600
rect 2590 6570 2650 6580
rect 2760 6600 2820 6610
rect 2760 6580 2770 6600
rect 2810 6580 2820 6600
rect 2760 6570 2820 6580
rect 2930 6600 2990 6610
rect 2930 6580 2940 6600
rect 2980 6580 2990 6600
rect 2930 6570 2990 6580
rect 3100 6600 3160 6610
rect 3100 6580 3110 6600
rect 3150 6580 3160 6600
rect 3100 6570 3160 6580
rect 3270 6600 3330 6610
rect 3500 6600 3560 6610
rect 3270 6580 3280 6600
rect 3320 6580 3510 6600
rect 3550 6580 3560 6600
rect 3270 6570 3330 6580
rect 3500 6570 3560 6580
rect 3500 6060 3560 6070
rect 3460 6040 3510 6060
rect 3550 6040 3560 6060
rect 1740 5560 1800 5570
rect 1740 5540 1750 5560
rect 1790 5540 1800 5560
rect 1910 5560 1970 5570
rect 1910 5540 1920 5560
rect 1960 5540 1970 5560
rect 2080 5560 2140 5570
rect 2080 5540 2090 5560
rect 2130 5540 2140 5560
rect 2250 5560 2310 5570
rect 2250 5540 2260 5560
rect 2300 5540 2310 5560
rect 2420 5560 2480 5570
rect 2420 5540 2430 5560
rect 2470 5540 2480 5560
rect 2590 5560 2650 5570
rect 2590 5540 2600 5560
rect 2640 5540 2650 5560
rect 2760 5560 2820 5570
rect 2760 5540 2770 5560
rect 2810 5540 2820 5560
rect 2930 5560 2990 5570
rect 2930 5540 2940 5560
rect 2980 5540 2990 5560
rect 3100 5560 3160 5570
rect 3100 5540 3110 5560
rect 3150 5540 3160 5560
rect 3270 5560 3330 5570
rect 3270 5540 3280 5560
rect 3320 5540 3330 5560
rect -10 5520 3330 5540
rect -10 5500 0 5520
rect 40 5500 50 5520
rect -10 5490 50 5500
rect 160 5500 170 5520
rect 210 5500 220 5520
rect 160 5490 220 5500
rect 330 5500 340 5520
rect 380 5500 390 5520
rect 330 5490 390 5500
rect 500 5500 510 5520
rect 550 5500 560 5520
rect 500 5490 560 5500
rect 670 5500 680 5520
rect 720 5500 730 5520
rect 670 5490 730 5500
rect 840 5500 850 5520
rect 890 5500 900 5520
rect 840 5490 900 5500
rect 1010 5500 1020 5520
rect 1060 5500 1070 5520
rect 1010 5490 1070 5500
rect 1180 5500 1190 5520
rect 1230 5500 1240 5520
rect 1180 5490 1240 5500
rect 1350 5500 1360 5520
rect 1400 5500 1410 5520
rect 1350 5490 1410 5500
rect 1520 5500 1530 5520
rect 1570 5500 1580 5520
rect 1520 5490 1580 5500
rect -120 5460 -80 5470
rect -120 5440 -110 5460
rect -90 5440 -80 5460
rect -120 5430 -80 5440
rect -110 5350 -90 5430
rect -10 5350 50 5360
rect 160 5350 220 5360
rect 330 5350 390 5360
rect 500 5350 560 5360
rect 670 5350 730 5360
rect 840 5350 900 5360
rect 1010 5350 1070 5360
rect 1180 5350 1240 5360
rect 1350 5350 1410 5360
rect 1520 5350 1580 5360
rect -110 5330 0 5350
rect 40 5330 170 5350
rect 210 5330 340 5350
rect 380 5330 510 5350
rect 550 5330 680 5350
rect 720 5330 850 5350
rect 890 5330 1020 5350
rect 1060 5330 1190 5350
rect 1230 5330 1360 5350
rect 1400 5330 1530 5350
rect 1570 5330 1580 5350
rect -10 5320 50 5330
rect 160 5320 220 5330
rect 330 5320 390 5330
rect 500 5320 560 5330
rect 670 5320 730 5330
rect 840 5320 900 5330
rect 1010 5320 1070 5330
rect 1180 5320 1240 5330
rect 1350 5320 1410 5330
rect 1520 5320 1580 5330
rect -230 5290 -190 5300
rect -160 5290 -60 5310
rect -230 5270 -220 5290
rect -200 5270 -190 5290
rect -230 5260 -190 5270
rect -220 5220 -200 5260
rect -80 5220 -60 5290
rect 50 5290 90 5300
rect 330 5290 370 5300
rect 610 5290 650 5300
rect 890 5290 930 5300
rect 1170 5290 1210 5300
rect 1520 5290 1540 5320
rect 50 5270 60 5290
rect 80 5270 340 5290
rect 360 5270 620 5290
rect 640 5270 900 5290
rect 920 5270 1180 5290
rect 1200 5270 1540 5290
rect 50 5260 90 5270
rect 330 5260 370 5270
rect 610 5260 650 5270
rect 890 5260 930 5270
rect 1170 5260 1210 5270
rect 60 5220 80 5260
rect 340 5220 360 5260
rect 620 5220 640 5260
rect 900 5220 920 5260
rect 1180 5220 1200 5260
rect 1520 5250 1540 5270
rect 1580 5290 1620 5300
rect 1580 5270 1590 5290
rect 1610 5270 1620 5290
rect 1580 5260 1620 5270
rect 1520 5240 1560 5250
rect 1520 5220 1530 5240
rect 1550 5220 1560 5240
rect -270 5210 -190 5220
rect -270 5170 -260 5210
rect -240 5170 -220 5210
rect -200 5170 -190 5210
rect -270 5160 -190 5170
rect -90 5210 -50 5220
rect -90 5170 -80 5210
rect -60 5170 -50 5210
rect -90 5160 -50 5170
rect 50 5210 90 5220
rect 50 5170 60 5210
rect 80 5170 90 5210
rect 50 5160 90 5170
rect 190 5210 230 5220
rect 190 5170 200 5210
rect 220 5170 230 5210
rect 190 5160 230 5170
rect 330 5210 370 5220
rect 330 5170 340 5210
rect 360 5170 370 5210
rect 330 5160 370 5170
rect 470 5210 510 5220
rect 470 5170 480 5210
rect 500 5170 510 5210
rect 470 5160 510 5170
rect 610 5210 650 5220
rect 610 5170 620 5210
rect 640 5170 650 5210
rect 610 5160 650 5170
rect 750 5210 790 5220
rect 750 5170 760 5210
rect 780 5170 790 5210
rect 750 5160 790 5170
rect 890 5210 930 5220
rect 890 5170 900 5210
rect 920 5170 930 5210
rect 890 5160 930 5170
rect 1030 5210 1070 5220
rect 1030 5170 1040 5210
rect 1060 5170 1070 5210
rect 1030 5160 1070 5170
rect 1170 5210 1210 5220
rect 1170 5170 1180 5210
rect 1200 5170 1210 5210
rect 1170 5160 1210 5170
rect 1310 5210 1350 5220
rect 1520 5210 1560 5220
rect 1310 5170 1320 5210
rect 1340 5180 1350 5210
rect 1340 5170 1560 5180
rect 1310 5160 1530 5170
rect -220 5100 -200 5160
rect -80 5140 -60 5160
rect 200 5140 220 5160
rect 480 5140 500 5160
rect 760 5140 780 5160
rect 1040 5140 1060 5160
rect 1320 5140 1340 5160
rect 1520 5150 1530 5160
rect 1550 5150 1560 5170
rect 1520 5140 1560 5150
rect -80 5120 1340 5140
rect 1380 5100 1420 5110
rect 1520 5100 1560 5110
rect -220 5080 1390 5100
rect 1410 5080 1530 5100
rect 1550 5080 1560 5100
rect -220 5020 -200 5080
rect 1380 5070 1420 5080
rect 1520 5070 1560 5080
rect -80 5040 1340 5060
rect -80 5020 -60 5040
rect 200 5020 220 5040
rect 480 5020 500 5040
rect 760 5020 780 5040
rect 1040 5020 1060 5040
rect 1320 5020 1340 5040
rect 1520 5030 1560 5040
rect 1520 5020 1530 5030
rect -270 5010 -190 5020
rect -270 4970 -260 5010
rect -240 4970 -220 5010
rect -200 4970 -190 5010
rect -270 4960 -190 4970
rect -90 5010 -50 5020
rect -90 4970 -80 5010
rect -60 4970 -50 5010
rect -90 4960 -50 4970
rect 50 5010 90 5020
rect 50 4970 60 5010
rect 80 4970 90 5010
rect 50 4960 90 4970
rect 190 5010 230 5020
rect 190 4970 200 5010
rect 220 4970 230 5010
rect 190 4960 230 4970
rect 330 5010 370 5020
rect 330 4970 340 5010
rect 360 4970 370 5010
rect 330 4960 370 4970
rect 470 5010 510 5020
rect 470 4970 480 5010
rect 500 4970 510 5010
rect 470 4960 510 4970
rect 610 5010 650 5020
rect 610 4970 620 5010
rect 640 4970 650 5010
rect 610 4960 650 4970
rect 750 5010 790 5020
rect 750 4970 760 5010
rect 780 4970 790 5010
rect 750 4960 790 4970
rect 890 5010 930 5020
rect 890 4970 900 5010
rect 920 4970 930 5010
rect 890 4960 930 4970
rect 1030 5010 1070 5020
rect 1030 4970 1040 5010
rect 1060 4970 1070 5010
rect 1030 4960 1070 4970
rect 1170 5010 1210 5020
rect 1170 4970 1180 5010
rect 1200 4970 1210 5010
rect 1170 4960 1210 4970
rect 1310 5010 1530 5020
rect 1550 5010 1560 5030
rect 1310 4970 1320 5010
rect 1340 5000 1560 5010
rect 1340 4970 1350 5000
rect 1310 4960 1350 4970
rect 1520 4960 1560 4970
rect -220 4920 -200 4960
rect -230 4910 -190 4920
rect -230 4890 -220 4910
rect -200 4890 -190 4910
rect -80 4890 -60 4960
rect 60 4920 80 4960
rect 340 4920 360 4960
rect 620 4920 640 4960
rect 900 4920 920 4960
rect 1180 4920 1200 4960
rect 1520 4940 1530 4960
rect 1550 4940 1560 4960
rect 1520 4930 1560 4940
rect -230 4880 -190 4890
rect -220 4690 -200 4880
rect -160 4870 -60 4890
rect 50 4910 90 4920
rect 330 4910 370 4920
rect 610 4910 650 4920
rect 890 4910 930 4920
rect 1170 4910 1210 4920
rect 1520 4910 1540 4930
rect 1590 4920 1610 5260
rect 50 4890 60 4910
rect 80 4890 340 4910
rect 360 4890 620 4910
rect 640 4890 900 4910
rect 920 4890 1180 4910
rect 1200 4890 1540 4910
rect 50 4880 90 4890
rect 330 4880 370 4890
rect 610 4880 650 4890
rect 890 4880 930 4890
rect 1170 4880 1210 4890
rect -240 4680 -180 4690
rect -240 4660 -230 4680
rect -190 4660 -180 4680
rect -240 4650 -180 4660
rect -240 4140 -180 4150
rect -160 4140 -140 4870
rect 1520 4860 1540 4890
rect 1580 4910 1620 4920
rect 1580 4890 1590 4910
rect 1610 4890 1620 4910
rect 1580 4880 1620 4890
rect -10 4850 50 4860
rect 160 4850 220 4860
rect 330 4850 390 4860
rect 500 4850 560 4860
rect 670 4850 730 4860
rect 840 4850 900 4860
rect 1010 4850 1070 4860
rect 1180 4850 1240 4860
rect 1350 4850 1410 4860
rect 1520 4850 1580 4860
rect -110 4830 0 4850
rect 40 4830 170 4850
rect 210 4830 340 4850
rect 380 4830 510 4850
rect 550 4830 680 4850
rect 720 4830 850 4850
rect 890 4830 1020 4850
rect 1060 4830 1190 4850
rect 1230 4830 1360 4850
rect 1400 4830 1530 4850
rect 1570 4830 1580 4850
rect -110 4750 -90 4830
rect -10 4820 50 4830
rect 160 4820 220 4830
rect 330 4820 390 4830
rect 500 4820 560 4830
rect 670 4820 730 4830
rect 840 4820 900 4830
rect 1010 4820 1070 4830
rect 1180 4820 1240 4830
rect 1350 4820 1410 4830
rect 1520 4820 1580 4830
rect -120 4740 -80 4750
rect -120 4720 -110 4740
rect -90 4720 -80 4740
rect -120 4710 -80 4720
rect -10 4680 50 4690
rect -10 4660 0 4680
rect 40 4660 50 4680
rect 160 4680 220 4690
rect 160 4660 170 4680
rect 210 4660 220 4680
rect 330 4680 390 4690
rect 330 4660 340 4680
rect 380 4660 390 4680
rect 500 4680 560 4690
rect 500 4660 510 4680
rect 550 4660 560 4680
rect 670 4680 730 4690
rect 670 4660 680 4680
rect 720 4660 730 4680
rect 840 4680 900 4690
rect 840 4660 850 4680
rect 890 4660 900 4680
rect 1010 4680 1070 4690
rect 1010 4660 1020 4680
rect 1060 4660 1070 4680
rect 1180 4680 1240 4690
rect 1180 4660 1190 4680
rect 1230 4660 1240 4680
rect 1350 4680 1410 4690
rect 1350 4660 1360 4680
rect 1400 4660 1410 4680
rect 1520 4680 1580 4690
rect 1520 4660 1530 4680
rect 1570 4660 1580 4680
rect 1650 4660 1670 5520
rect 1740 5500 1750 5520
rect 1790 5500 1800 5520
rect 1740 5490 1800 5500
rect 1910 5500 1920 5520
rect 1960 5500 1970 5520
rect 1910 5490 1970 5500
rect 2080 5500 2090 5520
rect 2130 5500 2140 5520
rect 2080 5490 2140 5500
rect 2250 5500 2260 5520
rect 2300 5500 2310 5520
rect 2250 5490 2310 5500
rect 2420 5500 2430 5520
rect 2470 5500 2480 5520
rect 2420 5490 2480 5500
rect 2590 5500 2600 5520
rect 2640 5500 2650 5520
rect 2590 5490 2650 5500
rect 2760 5500 2770 5520
rect 2810 5500 2820 5520
rect 2760 5490 2820 5500
rect 2930 5500 2940 5520
rect 2980 5500 2990 5520
rect 2930 5490 2990 5500
rect 3100 5500 3110 5520
rect 3150 5500 3160 5520
rect 3100 5490 3160 5500
rect 3270 5500 3280 5520
rect 3320 5500 3330 5520
rect 3270 5490 3330 5500
rect 3400 5460 3440 5470
rect 3400 5440 3410 5460
rect 3430 5440 3440 5460
rect 3400 5430 3440 5440
rect 1740 5350 1800 5360
rect 1910 5350 1970 5360
rect 2080 5350 2140 5360
rect 2250 5350 2310 5360
rect 2420 5350 2480 5360
rect 2590 5350 2650 5360
rect 2760 5350 2820 5360
rect 2930 5350 2990 5360
rect 3100 5350 3160 5360
rect 3270 5350 3330 5360
rect 3410 5350 3430 5430
rect 1740 5330 1750 5350
rect 1790 5330 1920 5350
rect 1960 5330 2090 5350
rect 2130 5330 2260 5350
rect 2300 5330 2430 5350
rect 2470 5330 2600 5350
rect 2640 5330 2770 5350
rect 2810 5330 2940 5350
rect 2980 5330 3110 5350
rect 3150 5330 3280 5350
rect 3320 5330 3430 5350
rect 1740 5320 1800 5330
rect 1910 5320 1970 5330
rect 2080 5320 2140 5330
rect 2250 5320 2310 5330
rect 2420 5320 2480 5330
rect 2590 5320 2650 5330
rect 2760 5320 2820 5330
rect 2930 5320 2990 5330
rect 3100 5320 3160 5330
rect 3270 5320 3330 5330
rect 1700 5290 1740 5300
rect 1700 5270 1710 5290
rect 1730 5270 1740 5290
rect 1700 5260 1740 5270
rect 1780 5290 1800 5320
rect 3460 5310 3480 6040
rect 3500 6030 3560 6040
rect 3500 5520 3560 5530
rect 3500 5500 3510 5520
rect 3550 5500 3560 5520
rect 3500 5490 3560 5500
rect 2110 5290 2150 5300
rect 2390 5290 2430 5300
rect 2670 5290 2710 5300
rect 2950 5290 2990 5300
rect 3230 5290 3270 5300
rect 1780 5270 2120 5290
rect 2140 5270 2400 5290
rect 2420 5270 2680 5290
rect 2700 5270 2960 5290
rect 2980 5270 3240 5290
rect 3260 5270 3270 5290
rect 1710 4920 1730 5260
rect 1780 5250 1800 5270
rect 2110 5260 2150 5270
rect 2390 5260 2430 5270
rect 2670 5260 2710 5270
rect 2950 5260 2990 5270
rect 3230 5260 3270 5270
rect 3380 5290 3480 5310
rect 3520 5300 3540 5490
rect 3510 5290 3550 5300
rect 1760 5240 1800 5250
rect 1760 5220 1770 5240
rect 1790 5220 1800 5240
rect 2120 5220 2140 5260
rect 2400 5220 2420 5260
rect 2680 5220 2700 5260
rect 2960 5220 2980 5260
rect 3240 5220 3260 5260
rect 3380 5220 3400 5290
rect 3510 5270 3520 5290
rect 3540 5270 3550 5290
rect 3510 5260 3550 5270
rect 3520 5220 3540 5260
rect 1760 5210 1800 5220
rect 1970 5210 2010 5220
rect 1970 5180 1980 5210
rect 1760 5170 1980 5180
rect 2000 5170 2010 5210
rect 1760 5150 1770 5170
rect 1790 5160 2010 5170
rect 2110 5210 2150 5220
rect 2110 5170 2120 5210
rect 2140 5170 2150 5210
rect 2110 5160 2150 5170
rect 2250 5210 2290 5220
rect 2250 5170 2260 5210
rect 2280 5170 2290 5210
rect 2250 5160 2290 5170
rect 2390 5210 2430 5220
rect 2390 5170 2400 5210
rect 2420 5170 2430 5210
rect 2390 5160 2430 5170
rect 2530 5210 2570 5220
rect 2530 5170 2540 5210
rect 2560 5170 2570 5210
rect 2530 5160 2570 5170
rect 2670 5210 2710 5220
rect 2670 5170 2680 5210
rect 2700 5170 2710 5210
rect 2670 5160 2710 5170
rect 2810 5210 2850 5220
rect 2810 5170 2820 5210
rect 2840 5170 2850 5210
rect 2810 5160 2850 5170
rect 2950 5210 2990 5220
rect 2950 5170 2960 5210
rect 2980 5170 2990 5210
rect 2950 5160 2990 5170
rect 3090 5210 3130 5220
rect 3090 5170 3100 5210
rect 3120 5170 3130 5210
rect 3090 5160 3130 5170
rect 3230 5210 3270 5220
rect 3230 5170 3240 5210
rect 3260 5170 3270 5210
rect 3230 5160 3270 5170
rect 3370 5210 3410 5220
rect 3370 5170 3380 5210
rect 3400 5170 3410 5210
rect 3370 5160 3410 5170
rect 3510 5210 3590 5220
rect 3510 5170 3520 5210
rect 3540 5170 3560 5210
rect 3580 5170 3590 5210
rect 3510 5160 3590 5170
rect 1790 5150 1800 5160
rect 1760 5140 1800 5150
rect 1980 5140 2000 5160
rect 2260 5140 2280 5160
rect 2540 5140 2560 5160
rect 2820 5140 2840 5160
rect 3100 5140 3120 5160
rect 3380 5140 3400 5160
rect 1980 5120 3400 5140
rect 1760 5100 1800 5110
rect 1900 5100 1940 5110
rect 3520 5100 3540 5160
rect 1760 5080 1770 5100
rect 1790 5080 1910 5100
rect 1930 5080 3540 5100
rect 1760 5070 1800 5080
rect 1900 5070 1940 5080
rect 1980 5040 3400 5060
rect 1760 5030 1800 5040
rect 1760 5010 1770 5030
rect 1790 5020 1800 5030
rect 1980 5020 2000 5040
rect 2260 5020 2280 5040
rect 2540 5020 2560 5040
rect 2820 5020 2840 5040
rect 3100 5020 3120 5040
rect 3380 5020 3400 5040
rect 3520 5020 3540 5080
rect 1790 5010 2010 5020
rect 1760 5000 1980 5010
rect 1970 4970 1980 5000
rect 2000 4970 2010 5010
rect 1760 4960 1800 4970
rect 1970 4960 2010 4970
rect 2110 5010 2150 5020
rect 2110 4970 2120 5010
rect 2140 4970 2150 5010
rect 2110 4960 2150 4970
rect 2250 5010 2290 5020
rect 2250 4970 2260 5010
rect 2280 4970 2290 5010
rect 2250 4960 2290 4970
rect 2390 5010 2430 5020
rect 2390 4970 2400 5010
rect 2420 4970 2430 5010
rect 2390 4960 2430 4970
rect 2530 5010 2570 5020
rect 2530 4970 2540 5010
rect 2560 4970 2570 5010
rect 2530 4960 2570 4970
rect 2670 5010 2710 5020
rect 2670 4970 2680 5010
rect 2700 4970 2710 5010
rect 2670 4960 2710 4970
rect 2810 5010 2850 5020
rect 2810 4970 2820 5010
rect 2840 4970 2850 5010
rect 2810 4960 2850 4970
rect 2950 5010 2990 5020
rect 2950 4970 2960 5010
rect 2980 4970 2990 5010
rect 2950 4960 2990 4970
rect 3090 5010 3130 5020
rect 3090 4970 3100 5010
rect 3120 4970 3130 5010
rect 3090 4960 3130 4970
rect 3230 5010 3270 5020
rect 3230 4970 3240 5010
rect 3260 4970 3270 5010
rect 3230 4960 3270 4970
rect 3370 5010 3410 5020
rect 3370 4970 3380 5010
rect 3400 4970 3410 5010
rect 3370 4960 3410 4970
rect 3510 5010 3590 5020
rect 3510 4970 3520 5010
rect 3540 4970 3560 5010
rect 3580 4970 3590 5010
rect 3510 4960 3590 4970
rect 1760 4940 1770 4960
rect 1790 4940 1800 4960
rect 1760 4930 1800 4940
rect 1700 4910 1740 4920
rect 1700 4890 1710 4910
rect 1730 4890 1740 4910
rect 1700 4880 1740 4890
rect 1780 4910 1800 4930
rect 2120 4920 2140 4960
rect 2400 4920 2420 4960
rect 2680 4920 2700 4960
rect 2960 4920 2980 4960
rect 3240 4920 3260 4960
rect 2110 4910 2150 4920
rect 2390 4910 2430 4920
rect 2670 4910 2710 4920
rect 2950 4910 2990 4920
rect 3230 4910 3270 4920
rect 1780 4890 2120 4910
rect 2140 4890 2400 4910
rect 2420 4890 2680 4910
rect 2700 4890 2960 4910
rect 2980 4890 3240 4910
rect 3260 4890 3270 4910
rect 1780 4860 1800 4890
rect 2110 4880 2150 4890
rect 2390 4880 2430 4890
rect 2670 4880 2710 4890
rect 2950 4880 2990 4890
rect 3230 4880 3270 4890
rect 3380 4890 3400 4960
rect 3520 4920 3540 4960
rect 3510 4910 3550 4920
rect 3510 4890 3520 4910
rect 3540 4890 3550 4910
rect 3380 4870 3480 4890
rect 3510 4880 3550 4890
rect 1740 4850 1800 4860
rect 1910 4850 1970 4860
rect 2080 4850 2140 4860
rect 2250 4850 2310 4860
rect 2420 4850 2480 4860
rect 2590 4850 2650 4860
rect 2760 4850 2820 4860
rect 2930 4850 2990 4860
rect 3100 4850 3160 4860
rect 3270 4850 3330 4860
rect 1740 4830 1750 4850
rect 1790 4830 1920 4850
rect 1960 4830 2090 4850
rect 2130 4830 2260 4850
rect 2300 4830 2430 4850
rect 2470 4830 2600 4850
rect 2640 4830 2770 4850
rect 2810 4830 2940 4850
rect 2980 4830 3110 4850
rect 3150 4830 3280 4850
rect 3320 4830 3430 4850
rect 1740 4820 1800 4830
rect 1910 4820 1970 4830
rect 2080 4820 2140 4830
rect 2250 4820 2310 4830
rect 2420 4820 2480 4830
rect 2590 4820 2650 4830
rect 2760 4820 2820 4830
rect 2930 4820 2990 4830
rect 3100 4820 3160 4830
rect 3270 4820 3330 4830
rect 3410 4750 3430 4830
rect 3400 4740 3440 4750
rect 3400 4720 3410 4740
rect 3430 4720 3440 4740
rect 3400 4710 3440 4720
rect 1740 4680 1800 4690
rect 1740 4660 1750 4680
rect 1790 4660 1800 4680
rect 1910 4680 1970 4690
rect 1910 4660 1920 4680
rect 1960 4660 1970 4680
rect 2080 4680 2140 4690
rect 2080 4660 2090 4680
rect 2130 4660 2140 4680
rect 2250 4680 2310 4690
rect 2250 4660 2260 4680
rect 2300 4660 2310 4680
rect 2420 4680 2480 4690
rect 2420 4660 2430 4680
rect 2470 4660 2480 4680
rect 2590 4680 2650 4690
rect 2590 4660 2600 4680
rect 2640 4660 2650 4680
rect 2760 4680 2820 4690
rect 2760 4660 2770 4680
rect 2810 4660 2820 4680
rect 2930 4680 2990 4690
rect 2930 4660 2940 4680
rect 2980 4660 2990 4680
rect 3100 4680 3160 4690
rect 3100 4660 3110 4680
rect 3150 4660 3160 4680
rect 3270 4680 3330 4690
rect 3270 4660 3280 4680
rect 3320 4660 3330 4680
rect -10 4640 3330 4660
rect -10 4620 0 4640
rect 40 4620 50 4640
rect -10 4610 50 4620
rect 160 4620 170 4640
rect 210 4620 220 4640
rect 160 4610 220 4620
rect 330 4620 340 4640
rect 380 4620 390 4640
rect 330 4610 390 4620
rect 500 4620 510 4640
rect 550 4620 560 4640
rect 500 4610 560 4620
rect 670 4620 680 4640
rect 720 4620 730 4640
rect 670 4610 730 4620
rect 840 4620 850 4640
rect 890 4620 900 4640
rect 840 4610 900 4620
rect 1010 4620 1020 4640
rect 1060 4620 1070 4640
rect 1010 4610 1070 4620
rect 1180 4620 1190 4640
rect 1230 4620 1240 4640
rect 1180 4610 1240 4620
rect 1350 4620 1360 4640
rect 1400 4620 1410 4640
rect 1350 4610 1410 4620
rect 1520 4620 1530 4640
rect 1570 4620 1580 4640
rect 1520 4610 1580 4620
rect -240 4120 -230 4140
rect -190 4120 -140 4140
rect -240 4110 -180 4120
rect -240 3600 -180 3610
rect -10 3600 50 3610
rect -240 3580 -230 3600
rect -190 3580 0 3600
rect 40 3580 50 3600
rect -240 3570 -180 3580
rect -10 3570 50 3580
rect 160 3600 220 3610
rect 160 3580 170 3600
rect 210 3580 220 3600
rect 160 3570 220 3580
rect 330 3600 390 3610
rect 330 3580 340 3600
rect 380 3580 390 3600
rect 330 3570 390 3580
rect 500 3600 560 3610
rect 500 3580 510 3600
rect 550 3580 560 3600
rect 500 3570 560 3580
rect 670 3600 730 3610
rect 670 3580 680 3600
rect 720 3580 730 3600
rect 670 3570 730 3580
rect 840 3600 900 3610
rect 840 3580 850 3600
rect 890 3580 900 3600
rect 840 3570 900 3580
rect 1010 3600 1070 3610
rect 1010 3580 1020 3600
rect 1060 3580 1070 3600
rect 1010 3570 1070 3580
rect 1180 3600 1240 3610
rect 1180 3580 1190 3600
rect 1230 3580 1240 3600
rect 1180 3570 1240 3580
rect 1350 3600 1410 3610
rect 1350 3580 1360 3600
rect 1400 3580 1410 3600
rect 1350 3570 1410 3580
rect 1520 3600 1580 3610
rect 1520 3580 1530 3600
rect 1570 3580 1580 3600
rect 1520 3570 1580 3580
rect -340 3540 -300 3550
rect -220 3540 -200 3570
rect -340 3520 -330 3540
rect -310 3520 -200 3540
rect -340 3510 -300 3520
rect -10 2560 50 2570
rect -90 2540 -50 2550
rect -10 2540 0 2560
rect 40 2540 50 2560
rect 160 2560 220 2570
rect 160 2540 170 2560
rect 210 2540 220 2560
rect 330 2560 390 2570
rect 330 2540 340 2560
rect 380 2540 390 2560
rect 500 2560 560 2570
rect 500 2540 510 2560
rect 550 2540 560 2560
rect 670 2560 730 2570
rect 670 2540 680 2560
rect 720 2540 730 2560
rect 840 2560 900 2570
rect 840 2540 850 2560
rect 890 2540 900 2560
rect 1010 2560 1070 2570
rect 1010 2540 1020 2560
rect 1060 2540 1070 2560
rect 1180 2560 1240 2570
rect 1180 2540 1190 2560
rect 1230 2540 1240 2560
rect 1350 2560 1410 2570
rect 1350 2540 1360 2560
rect 1400 2540 1410 2560
rect 1520 2560 1580 2570
rect 1520 2540 1530 2560
rect 1570 2540 1580 2560
rect 1650 2540 1670 4640
rect 1740 4620 1750 4640
rect 1790 4620 1800 4640
rect 1740 4610 1800 4620
rect 1910 4620 1920 4640
rect 1960 4620 1970 4640
rect 1910 4610 1970 4620
rect 2080 4620 2090 4640
rect 2130 4620 2140 4640
rect 2080 4610 2140 4620
rect 2250 4620 2260 4640
rect 2300 4620 2310 4640
rect 2250 4610 2310 4620
rect 2420 4620 2430 4640
rect 2470 4620 2480 4640
rect 2420 4610 2480 4620
rect 2590 4620 2600 4640
rect 2640 4620 2650 4640
rect 2590 4610 2650 4620
rect 2760 4620 2770 4640
rect 2810 4620 2820 4640
rect 2760 4610 2820 4620
rect 2930 4620 2940 4640
rect 2980 4620 2990 4640
rect 2930 4610 2990 4620
rect 3100 4620 3110 4640
rect 3150 4620 3160 4640
rect 3100 4610 3160 4620
rect 3270 4620 3280 4640
rect 3320 4620 3330 4640
rect 3270 4610 3330 4620
rect 3460 4140 3480 4870
rect 3520 4690 3540 4880
rect 3500 4680 3560 4690
rect 3500 4660 3510 4680
rect 3550 4660 3560 4680
rect 3500 4650 3560 4660
rect 3500 4140 3560 4150
rect 3460 4120 3510 4140
rect 3550 4120 3560 4140
rect 3500 4110 3560 4120
rect 1740 3600 1800 3610
rect 1740 3580 1750 3600
rect 1790 3580 1800 3600
rect 1740 3570 1800 3580
rect 1910 3600 1970 3610
rect 1910 3580 1920 3600
rect 1960 3580 1970 3600
rect 1910 3570 1970 3580
rect 2080 3600 2140 3610
rect 2080 3580 2090 3600
rect 2130 3580 2140 3600
rect 2080 3570 2140 3580
rect 2250 3600 2310 3610
rect 2250 3580 2260 3600
rect 2300 3580 2310 3600
rect 2250 3570 2310 3580
rect 2420 3600 2480 3610
rect 2420 3580 2430 3600
rect 2470 3580 2480 3600
rect 2420 3570 2480 3580
rect 2590 3600 2650 3610
rect 2590 3580 2600 3600
rect 2640 3580 2650 3600
rect 2590 3570 2650 3580
rect 2760 3600 2820 3610
rect 2760 3580 2770 3600
rect 2810 3580 2820 3600
rect 2760 3570 2820 3580
rect 2930 3600 2990 3610
rect 2930 3580 2940 3600
rect 2980 3580 2990 3600
rect 2930 3570 2990 3580
rect 3100 3600 3160 3610
rect 3100 3580 3110 3600
rect 3150 3580 3160 3600
rect 3100 3570 3160 3580
rect 3270 3600 3330 3610
rect 3500 3600 3560 3610
rect 3270 3580 3280 3600
rect 3320 3580 3510 3600
rect 3550 3580 3560 3600
rect 3270 3570 3330 3580
rect 3500 3570 3560 3580
rect 3520 3540 3540 3570
rect 3630 3550 3650 6630
rect 3620 3540 3660 3550
rect 3520 3520 3630 3540
rect 3650 3520 3660 3540
rect 3620 3510 3660 3520
rect 1740 2560 1800 2570
rect 1740 2540 1750 2560
rect 1790 2540 1800 2560
rect 1910 2560 1970 2570
rect 1910 2540 1920 2560
rect 1960 2540 1970 2560
rect 2080 2560 2140 2570
rect 2080 2540 2090 2560
rect 2130 2540 2140 2560
rect 2250 2560 2310 2570
rect 2250 2540 2260 2560
rect 2300 2540 2310 2560
rect 2420 2560 2480 2570
rect 2420 2540 2430 2560
rect 2470 2540 2480 2560
rect 2590 2560 2650 2570
rect 2590 2540 2600 2560
rect 2640 2540 2650 2560
rect 2760 2560 2820 2570
rect 2760 2540 2770 2560
rect 2810 2540 2820 2560
rect 2930 2560 2990 2570
rect 2930 2540 2940 2560
rect 2980 2540 2990 2560
rect 3100 2560 3160 2570
rect 3100 2540 3110 2560
rect 3150 2540 3160 2560
rect 3270 2560 3330 2570
rect 3270 2540 3280 2560
rect 3320 2540 3330 2560
rect 3370 2540 3410 2550
rect -90 2520 -80 2540
rect -60 2520 3380 2540
rect 3400 2520 3410 2540
rect -90 2510 -50 2520
rect -10 2500 0 2520
rect 40 2500 50 2520
rect 160 2500 170 2520
rect 210 2500 220 2520
rect 330 2500 340 2520
rect 380 2500 390 2520
rect 500 2500 510 2520
rect 550 2500 560 2520
rect 670 2500 680 2520
rect 720 2500 730 2520
rect 840 2500 850 2520
rect 890 2500 900 2520
rect 1010 2500 1020 2520
rect 1060 2500 1070 2520
rect 1180 2500 1190 2520
rect 1230 2500 1240 2520
rect 1350 2500 1360 2520
rect 1400 2500 1410 2520
rect 1520 2500 1530 2520
rect 1570 2500 1580 2520
rect 1740 2500 1750 2520
rect 1790 2500 1800 2520
rect 1910 2500 1920 2520
rect 1960 2500 1970 2520
rect 2080 2500 2090 2520
rect 2130 2500 2140 2520
rect 2250 2500 2260 2520
rect 2300 2500 2310 2520
rect 2420 2500 2430 2520
rect 2470 2500 2480 2520
rect 2590 2500 2600 2520
rect 2640 2500 2650 2520
rect 2760 2500 2770 2520
rect 2810 2500 2820 2520
rect 2930 2500 2940 2520
rect 2980 2500 2990 2520
rect 3100 2500 3110 2520
rect 3150 2500 3160 2520
rect 3270 2500 3280 2520
rect 3320 2500 3330 2520
rect 3370 2510 3410 2520
<< labels >>
rlabel locali -90 7650 -90 7650 7 VN
port 1 w
rlabel locali -220 5090 -220 5090 7 VP
port 2 w
rlabel locali -340 6650 -340 6650 7 Vc
port 3 w
rlabel locali 1720 5300 1720 5300 1 Vbn
port 4 n
rlabel locali 1800 5230 1800 5230 3 Vbg
rlabel locali 1780 5180 1780 5180 1 Vdssat
<< end >>
