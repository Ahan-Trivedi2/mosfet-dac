* SPICE3 file created from pcbc.ext - technology: sky130A


* Top level circuit pcbc

X0 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X1 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X2 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X3 a_8360_6840# a_8320_6920# w_8320_5720# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X4 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X5 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X6 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X7 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X8 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X9 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X10 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X11 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X12 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X13 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X14 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X15 a_8360_6840# a_8320_6920# w_8320_5720# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X16 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X17 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X18 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X19 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X20 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X21 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X22 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X23 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X24 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X25 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X26 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X27 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X28 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X29 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X30 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X31 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X32 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X33 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X34 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X35 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X36 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X37 w_8320_5720# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X38 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X39 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X40 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X41 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X42 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X43 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X44 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X45 a_8300_5640# a_8300_5640# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X46 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X47 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X48 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X49 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X50 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X51 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X52 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X53 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X54 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X55 a_8300_5640# a_8300_5640# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X56 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X57 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X58 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X59 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X60 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X61 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X62 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X63 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X64 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X65 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X66 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X67 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X68 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X69 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X70 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X71 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X72 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X73 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X74 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X75 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X76 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X77 a_8360_6840# a_8300_5640# a_8300_5640# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X78 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X79 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X80 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X81 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X82 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X83 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X84 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X85 w_8320_5720# w_8320_5720# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X86 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X87 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X88 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X89 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X90 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X91 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X92 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X93 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X94 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X95 w_8320_5720# w_8320_5720# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X96 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X97 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X98 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X99 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X100 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X101 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X102 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X103 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X104 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X105 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X106 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X107 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X108 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X109 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X110 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X111 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X112 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X113 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X114 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X115 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X116 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X117 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X118 a_8360_6840# w_8320_5720# w_8320_5720# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X119 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X120 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X121 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X122 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X123 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X124 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X125 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X126 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X127 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X128 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X129 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X130 w_8320_5720# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X131 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X132 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X133 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X134 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X135 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X136 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X137 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X138 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X139 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X140 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X141 a_8360_6840# w_8320_5720# w_8320_5720# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X142 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X143 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X144 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X145 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X146 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X147 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X148 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X149 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X150 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X151 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X152 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X153 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X154 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X155 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X156 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X157 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X158 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X159 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X160 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X161 a_8800_5440# a_8880_5840# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X162 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X163 a_8300_5640# a_8800_5440# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X164 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X165 a_8800_5440# a_8800_5440# a_8300_5640# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X166 a_8360_6840# a_8300_5640# a_8300_5640# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X167 a_8320_6920# a_8320_6920# a_8360_6840# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X168 a_8360_6840# a_8320_6920# a_8320_6920# w_8320_5720# sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X169 a_8300_5640# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X170 a_8800_5440# a_8880_5840# a_8320_6920# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X171 a_8320_6920# a_8880_5840# a_8800_5440# a_8800_5440# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
.end

