* SPICE3 file created from ncbc.ext - technology: sky130A

X0 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X1 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X2 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X3 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X4 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X5 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X6 Vdssat Vc Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X7 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X8 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X9 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X10 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X11 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X12 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X13 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X14 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X15 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X16 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X17 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X18 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X19 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X20 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X21 Vc Vc Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X22 Vdssat VN VN VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.56 ps=4.4 w=1 l=1
X23 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X24 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X25 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X26 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X27 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X28 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X29 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X30 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X31 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X32 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X33 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X34 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X35 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X36 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X37 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X38 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X39 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X40 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X41 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X42 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X43 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X44 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X45 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X46 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X47 VN Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X48 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X49 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X50 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.5 ps=3.6 w=1 l=1
X51 VN VN Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.56 pd=4.4 as=0.2 ps=1.4 w=1 l=1
X52 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X53 Vdssat VN VN VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.56 ps=4.4 w=1 l=1
X54 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X55 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X56 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X57 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X58 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X59 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X60 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X61 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X62 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X63 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X64 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X65 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X66 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X67 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X68 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X69 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X70 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X71 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X72 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3.6 as=0.5 ps=3.6 w=1 l=1
X73 Vdssat Vc Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X74 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X75 Vdssat Vbg VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X76 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X77 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X78 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X79 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X80 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X81 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X82 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X83 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.5 ps=3.6 w=1 l=1
X84 VN VN Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.56 pd=4.4 as=0.2 ps=1.4 w=1 l=1
X85 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X86 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X87 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X88 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X89 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X90 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X91 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X92 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3.6 as=0.2 ps=1.4 w=1 l=1
X93 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X94 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X95 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X96 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X97 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X98 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X99 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X100 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X101 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X102 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X103 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X104 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X105 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X106 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X107 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X108 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X109 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X110 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X111 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3.6 as=0.5 ps=3.6 w=1 l=1
X112 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X113 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X114 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X115 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X116 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X117 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3.6 as=0.5 ps=3.6 w=1 l=1
X118 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X119 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X120 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X121 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X122 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X123 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X124 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X125 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X126 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X127 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X128 VN Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X129 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X130 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3.6 as=0.2 ps=1.4 w=1 l=1
X131 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X132 Vc Vc Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X133 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X134 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X135 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X136 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X137 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X138 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X139 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X140 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X141 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X142 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X143 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X144 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X145 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X146 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X147 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X148 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X149 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3.6 as=0.5 ps=3.6 w=1 l=1
X150 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X151 Vdssat Vbg VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X152 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X153 Vdssat Vbg Vbg VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X154 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X155 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X156 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X157 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X158 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X159 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X160 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X161 Vbg Vbg Vdssat VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X162 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X163 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X164 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X165 VP Vbp Vc VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X166 Vbg Vbp VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X167 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X168 VP Vbp Vbg VP sky130_fd_pr__pfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X169 VP VP Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X170 Vc VP VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X171 Vc Vbp VP VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
.end

