magic
tech sky130A
timestamp 1762025964
<< nwell >>
rect -150 -160 325 200
rect 2715 -160 3190 200
<< nmos >>
rect 415 55 915 255
rect 965 55 1465 255
rect 1515 55 2015 255
rect 2065 55 2565 255
rect 415 -365 915 -165
rect 965 -365 1465 -165
rect 1515 -365 2015 -165
rect 2065 -365 2565 -165
<< pmos >>
rect 5 80 105 180
rect 155 80 255 180
rect 2870 80 2970 180
rect 3020 80 3120 180
rect 5 -140 105 -40
rect 155 -140 255 -40
rect 2870 -140 2970 -40
rect 3020 -140 3120 -40
<< ndiff >>
rect 365 240 415 255
rect 365 70 380 240
rect 400 70 415 240
rect 365 55 415 70
rect 915 240 965 255
rect 915 70 930 240
rect 950 70 965 240
rect 915 55 965 70
rect 1465 240 1515 255
rect 1465 70 1480 240
rect 1500 70 1515 240
rect 1465 55 1515 70
rect 2015 240 2065 255
rect 2015 70 2030 240
rect 2050 70 2065 240
rect 2015 55 2065 70
rect 2565 240 2615 255
rect 2565 70 2580 240
rect 2600 70 2615 240
rect 2565 55 2615 70
rect 365 -180 415 -165
rect 365 -350 380 -180
rect 400 -350 415 -180
rect 365 -365 415 -350
rect 915 -180 965 -165
rect 915 -350 930 -180
rect 950 -350 965 -180
rect 915 -365 965 -350
rect 1465 -180 1515 -165
rect 1465 -350 1480 -180
rect 1500 -350 1515 -180
rect 1465 -365 1515 -350
rect 2015 -180 2065 -165
rect 2015 -350 2030 -180
rect 2050 -350 2065 -180
rect 2015 -365 2065 -350
rect 2565 -180 2615 -165
rect 2565 -350 2580 -180
rect 2600 -350 2615 -180
rect 2565 -365 2615 -350
<< pdiff >>
rect -45 165 5 180
rect -45 95 -30 165
rect -10 95 5 165
rect -45 80 5 95
rect 105 165 155 180
rect 105 95 120 165
rect 140 95 155 165
rect 105 80 155 95
rect 255 165 305 180
rect 255 95 270 165
rect 290 95 305 165
rect 255 80 305 95
rect 2820 165 2870 180
rect 2820 95 2835 165
rect 2855 95 2870 165
rect 2820 80 2870 95
rect 2970 165 3020 180
rect 2970 95 2985 165
rect 3005 95 3020 165
rect 2970 80 3020 95
rect 3120 165 3170 180
rect 3120 95 3135 165
rect 3155 95 3170 165
rect 3120 80 3170 95
rect -45 -55 5 -40
rect -45 -125 -30 -55
rect -10 -125 5 -55
rect -45 -140 5 -125
rect 105 -55 155 -40
rect 105 -125 120 -55
rect 140 -125 155 -55
rect 105 -140 155 -125
rect 255 -55 305 -40
rect 255 -125 270 -55
rect 290 -125 305 -55
rect 255 -140 305 -125
rect 2820 -55 2870 -40
rect 2820 -125 2835 -55
rect 2855 -125 2870 -55
rect 2820 -140 2870 -125
rect 2970 -55 3020 -40
rect 2970 -125 2985 -55
rect 3005 -125 3020 -55
rect 2970 -140 3020 -125
rect 3120 -55 3170 -40
rect 3120 -125 3135 -55
rect 3155 -125 3170 -55
rect 3120 -140 3170 -125
<< ndiffc >>
rect 380 70 400 240
rect 930 70 950 240
rect 1480 70 1500 240
rect 2030 70 2050 240
rect 2580 70 2600 240
rect 380 -350 400 -180
rect 930 -350 950 -180
rect 1480 -350 1500 -180
rect 2030 -350 2050 -180
rect 2580 -350 2600 -180
<< pdiffc >>
rect -30 95 -10 165
rect 120 95 140 165
rect 270 95 290 165
rect 2835 95 2855 165
rect 2985 95 3005 165
rect 3135 95 3155 165
rect -30 -125 -10 -55
rect 120 -125 140 -55
rect 270 -125 290 -55
rect 2835 -125 2855 -55
rect 2985 -125 3005 -55
rect 3135 -125 3155 -55
<< psubdiff >>
rect 1530 -20 1580 -5
rect 1530 -90 1545 -20
rect 1565 -90 1580 -20
rect 1530 -105 1580 -90
<< nsubdiff >>
rect -130 -55 -80 -40
rect -130 -125 -115 -55
rect -95 -125 -80 -55
rect -130 -140 -80 -125
rect 2735 -55 2785 -40
rect 2735 -125 2750 -55
rect 2770 -125 2785 -55
rect 2735 -140 2785 -125
<< psubdiffcont >>
rect 1545 -90 1565 -20
<< nsubdiffcont >>
rect -115 -125 -95 -55
rect 2750 -125 2770 -55
<< poly >>
rect 415 255 915 270
rect 965 255 1465 270
rect 1515 255 2015 270
rect 2065 255 2565 270
rect 5 180 105 195
rect 155 180 255 195
rect 5 65 105 80
rect 155 65 255 80
rect 2870 180 2970 195
rect 3020 180 3120 195
rect 2870 65 2970 80
rect 3020 65 3120 80
rect 415 40 915 55
rect 965 40 1465 55
rect 1515 40 2015 55
rect 2065 40 2565 55
rect 5 -40 105 -25
rect 155 -40 255 -25
rect 2870 -40 2970 -25
rect 3020 -40 3120 -25
rect 5 -155 105 -140
rect 155 -155 255 -140
rect 415 -165 915 -150
rect 965 -165 1465 -150
rect 1515 -165 2015 -150
rect 2065 -165 2565 -150
rect 2870 -155 2970 -140
rect 3020 -155 3120 -140
rect 415 -380 915 -365
rect 965 -380 1465 -365
rect 1515 -380 2015 -365
rect 2065 -380 2565 -365
<< locali >>
rect 370 240 410 250
rect -40 165 0 175
rect -40 95 -30 165
rect -10 95 0 165
rect -40 85 0 95
rect 110 165 150 175
rect 110 95 120 165
rect 140 95 150 165
rect 110 85 150 95
rect 260 165 300 175
rect 260 95 270 165
rect 290 95 300 165
rect 260 85 300 95
rect 370 70 380 240
rect 400 70 410 240
rect 370 60 410 70
rect 920 240 960 250
rect 920 70 930 240
rect 950 70 960 240
rect 920 60 960 70
rect 1470 240 1510 250
rect 1470 70 1480 240
rect 1500 70 1510 240
rect 1470 60 1510 70
rect 2020 240 2060 250
rect 2020 70 2030 240
rect 2050 70 2060 240
rect 2020 60 2060 70
rect 2570 240 2610 250
rect 2570 70 2580 240
rect 2600 70 2610 240
rect 2825 165 2865 175
rect 2825 95 2835 165
rect 2855 95 2865 165
rect 2825 85 2865 95
rect 2975 165 3015 175
rect 2975 95 2985 165
rect 3005 95 3015 165
rect 2975 85 3015 95
rect 3125 165 3165 175
rect 3125 95 3135 165
rect 3155 95 3165 165
rect 3125 85 3165 95
rect 2570 60 2610 70
rect 1535 -20 1575 -10
rect -125 -55 -85 -45
rect -125 -125 -115 -55
rect -95 -125 -85 -55
rect -125 -135 -85 -125
rect -40 -55 0 -45
rect -40 -125 -30 -55
rect -10 -125 0 -55
rect -40 -135 0 -125
rect 110 -55 150 -45
rect 110 -125 120 -55
rect 140 -125 150 -55
rect 110 -135 150 -125
rect 260 -55 300 -45
rect 260 -125 270 -55
rect 290 -125 300 -55
rect 1535 -90 1545 -20
rect 1565 -90 1575 -20
rect 1535 -100 1575 -90
rect 2740 -55 2780 -45
rect 260 -135 300 -125
rect 2740 -125 2750 -55
rect 2770 -125 2780 -55
rect 2740 -135 2780 -125
rect 2825 -55 2865 -45
rect 2825 -125 2835 -55
rect 2855 -125 2865 -55
rect 2825 -135 2865 -125
rect 2975 -55 3015 -45
rect 2975 -125 2985 -55
rect 3005 -125 3015 -55
rect 2975 -135 3015 -125
rect 3125 -55 3165 -45
rect 3125 -125 3135 -55
rect 3155 -125 3165 -55
rect 3125 -135 3165 -125
rect 370 -180 410 -170
rect 370 -350 380 -180
rect 400 -350 410 -180
rect 370 -360 410 -350
rect 920 -180 960 -170
rect 920 -350 930 -180
rect 950 -350 960 -180
rect 920 -360 960 -350
rect 1470 -180 1510 -170
rect 1470 -350 1480 -180
rect 1500 -350 1510 -180
rect 1470 -360 1510 -350
rect 2020 -180 2060 -170
rect 2020 -350 2030 -180
rect 2050 -350 2060 -180
rect 2020 -360 2060 -350
rect 2570 -180 2610 -170
rect 2570 -350 2580 -180
rect 2600 -350 2610 -180
rect 2570 -360 2610 -350
<< end >>
