magic
tech sky130A
timestamp 1762208113
<< nwell >>
rect -100 1080 1200 1090
rect -1810 570 2910 1080
rect -1810 30 -620 570
rect 1720 30 2910 570
<< nmos >>
rect -540 320 -40 520
rect 0 320 500 520
rect 600 320 1100 520
rect 1140 320 1640 520
rect -540 50 -40 250
rect 0 50 500 250
rect 600 50 1100 250
rect 1140 50 1640 250
<< pmos >>
rect -1720 860 -1220 1060
rect -1180 860 -680 1060
rect -640 860 -140 1060
rect -100 860 400 1060
rect -1720 590 -1220 790
rect -1180 590 -680 790
rect -640 590 -140 790
rect -100 590 400 790
rect 700 860 1200 1060
rect 1240 860 1740 1060
rect 1780 860 2280 1060
rect 2320 860 2820 1060
rect 700 590 1200 790
rect 1240 590 1740 790
rect 1780 590 2280 790
rect 2320 590 2820 790
rect -1720 320 -1220 520
rect -1180 320 -680 520
rect 1780 320 2280 520
rect 2320 320 2820 520
rect -1720 50 -1220 250
rect -1180 50 -680 250
rect 1780 50 2280 250
rect 2320 50 2820 250
<< ndiff >>
rect -580 430 -540 520
rect -580 410 -570 430
rect -550 410 -540 430
rect -580 320 -540 410
rect -40 320 0 520
rect 500 380 600 520
rect 500 360 540 380
rect 560 360 600 380
rect 500 320 600 360
rect 1100 320 1140 520
rect 1640 430 1680 520
rect 1640 410 1650 430
rect 1670 410 1680 430
rect 1640 320 1680 410
rect -570 250 -550 320
rect -30 250 -10 320
rect 510 250 530 320
rect 570 250 590 320
rect 1110 250 1130 320
rect 1650 250 1670 320
rect -580 160 -540 250
rect -580 140 -570 160
rect -550 140 -540 160
rect -580 50 -540 140
rect -40 50 0 250
rect 500 160 600 250
rect 500 140 540 160
rect 560 140 600 160
rect 500 50 600 140
rect 1100 50 1140 250
rect 1640 160 1680 250
rect 1640 140 1650 160
rect 1670 140 1680 160
rect 1640 50 1680 140
<< pdiff >>
rect -1790 970 -1720 1060
rect -1790 950 -1750 970
rect -1730 950 -1720 970
rect -1790 860 -1720 950
rect -1220 970 -1180 1060
rect -1220 950 -1210 970
rect -1190 950 -1180 970
rect -1220 860 -1180 950
rect -680 860 -640 1060
rect -140 970 -100 1060
rect -140 950 -130 970
rect -110 950 -100 970
rect -140 860 -100 950
rect 400 970 470 1060
rect 400 950 410 970
rect 430 950 470 970
rect 630 970 700 1060
rect 400 860 470 950
rect -1750 790 -1730 860
rect -1210 790 -1190 860
rect -670 790 -650 860
rect -130 790 -110 860
rect 410 790 430 860
rect -1790 700 -1720 790
rect -1790 680 -1750 700
rect -1730 680 -1720 700
rect -1790 590 -1720 680
rect -1220 700 -1180 790
rect -1220 680 -1210 700
rect -1190 680 -1180 700
rect -1220 590 -1180 680
rect -680 590 -640 790
rect -140 700 -100 790
rect -140 680 -130 700
rect -110 680 -100 700
rect -140 590 -100 680
rect 400 700 470 790
rect 400 680 410 700
rect 430 680 470 700
rect 400 590 470 680
rect 630 950 670 970
rect 690 950 700 970
rect 630 860 700 950
rect 1200 970 1240 1060
rect 1200 950 1210 970
rect 1230 950 1240 970
rect 1200 860 1240 950
rect 1740 860 1780 1060
rect 2280 970 2320 1060
rect 2280 950 2290 970
rect 2310 950 2320 970
rect 2280 860 2320 950
rect 2820 970 2890 1060
rect 2820 950 2830 970
rect 2850 950 2890 970
rect 2820 860 2890 950
rect 670 790 690 860
rect 1210 790 1230 860
rect 1750 790 1770 860
rect 2290 790 2310 860
rect 2830 790 2850 860
rect 630 700 700 790
rect 630 680 670 700
rect 690 680 700 700
rect 630 590 700 680
rect 1200 700 1240 790
rect 1200 680 1210 700
rect 1230 680 1240 700
rect 1200 590 1240 680
rect 1740 590 1780 790
rect 2280 700 2320 790
rect 2280 680 2290 700
rect 2310 680 2320 700
rect 2280 590 2320 680
rect 2820 700 2890 790
rect 2820 680 2830 700
rect 2850 680 2890 700
rect 2820 590 2890 680
rect -1790 430 -1720 520
rect -1790 410 -1750 430
rect -1730 410 -1720 430
rect -1790 320 -1720 410
rect -1220 430 -1180 520
rect -1220 410 -1210 430
rect -1190 410 -1180 430
rect -1220 320 -1180 410
rect -680 430 -640 520
rect -680 410 -670 430
rect -650 410 -640 430
rect -680 320 -640 410
rect 1740 430 1780 520
rect 1740 410 1750 430
rect 1770 410 1780 430
rect 1740 320 1780 410
rect 2280 430 2320 520
rect 2280 410 2290 430
rect 2310 410 2320 430
rect 2280 320 2320 410
rect 2820 430 2890 520
rect 2820 410 2830 430
rect 2850 410 2890 430
rect 2820 320 2890 410
rect -1750 250 -1730 320
rect -1210 250 -1190 320
rect -670 250 -650 320
rect 1750 250 1770 320
rect 2290 250 2310 320
rect 2830 250 2850 320
rect -1790 160 -1720 250
rect -1790 140 -1750 160
rect -1730 140 -1720 160
rect -1790 50 -1720 140
rect -1220 160 -1180 250
rect -1220 140 -1210 160
rect -1190 140 -1180 160
rect -1220 50 -1180 140
rect -680 160 -640 250
rect -680 140 -670 160
rect -650 140 -640 160
rect -680 50 -640 140
rect 1740 160 1780 250
rect 1740 140 1750 160
rect 1770 140 1780 160
rect 1740 50 1780 140
rect 2280 160 2320 250
rect 2280 140 2290 160
rect 2310 140 2320 160
rect 2280 50 2320 140
rect 2820 160 2890 250
rect 2820 140 2830 160
rect 2850 140 2890 160
rect 2820 50 2890 140
<< ndiffc >>
rect -570 410 -550 430
rect 540 360 560 380
rect 1650 410 1670 430
rect -570 140 -550 160
rect 540 140 560 160
rect 1650 140 1670 160
<< pdiffc >>
rect -1750 950 -1730 970
rect -1210 950 -1190 970
rect -130 950 -110 970
rect 410 950 430 970
rect -1750 680 -1730 700
rect -1210 680 -1190 700
rect -130 680 -110 700
rect 410 680 430 700
rect 670 950 690 970
rect 1210 950 1230 970
rect 2290 950 2310 970
rect 2830 950 2850 970
rect 670 680 690 700
rect 1210 680 1230 700
rect 2290 680 2310 700
rect 2830 680 2850 700
rect -1750 410 -1730 430
rect -1210 410 -1190 430
rect -670 410 -650 430
rect 1750 410 1770 430
rect 2290 410 2310 430
rect 2830 410 2850 430
rect -1750 140 -1730 160
rect -1210 140 -1190 160
rect -670 140 -650 160
rect 1750 140 1770 160
rect 2290 140 2310 160
rect 2830 140 2850 160
<< psubdiff >>
rect 530 300 570 320
rect 530 270 540 300
rect 560 270 570 300
rect 530 250 570 270
<< nsubdiff >>
rect -1790 840 -1750 860
rect -1790 810 -1780 840
rect -1760 810 -1750 840
rect -1790 790 -1750 810
rect 430 840 470 860
rect 430 810 440 840
rect 460 810 470 840
rect 430 790 470 810
rect 630 840 670 860
rect 630 810 640 840
rect 660 810 670 840
rect 630 790 670 810
rect 2850 840 2890 860
rect 2850 810 2860 840
rect 2880 810 2890 840
rect 2850 790 2890 810
rect -1790 300 -1750 320
rect -1790 270 -1780 300
rect -1760 270 -1750 300
rect -1790 250 -1750 270
rect 2850 300 2890 320
rect 2850 270 2860 300
rect 2880 270 2890 300
rect 2850 250 2890 270
<< psubdiffcont >>
rect 540 270 560 300
<< nsubdiffcont >>
rect -1780 810 -1760 840
rect 440 810 460 840
rect 640 810 660 840
rect 2860 810 2880 840
rect -1780 270 -1760 300
rect 2860 270 2880 300
<< poly >>
rect -1260 1110 -1220 1120
rect -1260 1090 -1250 1110
rect -1230 1090 -1220 1110
rect -1260 1080 -1220 1090
rect -180 1110 -140 1120
rect -180 1090 -170 1110
rect -150 1090 -140 1110
rect 1240 1110 1280 1120
rect 1240 1090 1250 1110
rect 1270 1090 1280 1110
rect -180 1080 -140 1090
rect -1720 1060 -1220 1080
rect -1180 1060 -680 1080
rect -640 1060 -140 1080
rect -100 1070 1200 1090
rect -100 1060 400 1070
rect 530 990 570 1070
rect 700 1060 1200 1070
rect 1240 1080 1280 1090
rect 2320 1110 2360 1120
rect 2320 1090 2330 1110
rect 2350 1090 2360 1110
rect 2320 1080 2360 1090
rect 1240 1060 1740 1080
rect 1780 1060 2280 1080
rect 2320 1060 2820 1080
rect 530 970 540 990
rect 560 970 570 990
rect 530 960 570 970
rect -1720 840 -1220 860
rect -1690 810 -1650 840
rect -1590 810 -1550 840
rect -1490 810 -1450 840
rect -1390 810 -1350 840
rect -1290 810 -1250 840
rect -1720 790 -1220 810
rect -1180 840 -680 860
rect -1150 810 -1110 840
rect -1050 810 -1010 840
rect -950 810 -910 840
rect -850 810 -810 840
rect -750 810 -710 840
rect -1180 790 -680 810
rect -640 840 -140 860
rect -610 810 -570 840
rect -510 810 -470 840
rect -410 810 -370 840
rect -310 810 -270 840
rect -210 810 -170 840
rect -640 790 -140 810
rect -100 840 400 860
rect -70 810 -30 840
rect 30 810 70 840
rect 130 810 170 840
rect 230 810 270 840
rect 330 810 370 840
rect -100 790 400 810
rect 700 840 1200 860
rect 730 810 770 840
rect 830 810 870 840
rect 930 810 970 840
rect 1030 810 1070 840
rect 1130 810 1170 840
rect 700 790 1200 810
rect 1240 840 1740 860
rect 1270 810 1310 840
rect 1370 810 1410 840
rect 1470 810 1510 840
rect 1570 810 1610 840
rect 1670 810 1710 840
rect 1240 790 1740 810
rect 1780 840 2280 860
rect 1810 810 1850 840
rect 1910 810 1950 840
rect 2010 810 2050 840
rect 2110 810 2150 840
rect 2210 810 2250 840
rect 1780 790 2280 810
rect 2320 840 2820 860
rect 2350 810 2390 840
rect 2450 810 2490 840
rect 2550 810 2590 840
rect 2650 810 2690 840
rect 2750 810 2790 840
rect 2320 790 2820 810
rect -1720 570 -1220 590
rect -1180 570 -680 590
rect -640 570 -140 590
rect -100 570 400 590
rect 700 570 1200 590
rect 1240 570 1740 590
rect 1780 570 2280 590
rect 2320 570 2820 590
rect -1150 540 -1110 570
rect -1050 540 -1010 570
rect -950 540 -910 570
rect -850 540 -810 570
rect -750 540 -710 570
rect 1810 540 1850 570
rect 1910 540 1950 570
rect 2010 540 2050 570
rect 2110 540 2150 570
rect 2210 540 2250 570
rect -1720 520 -1220 540
rect -1180 520 -680 540
rect -540 520 -40 540
rect 0 520 500 540
rect 600 520 1100 540
rect 1140 520 1640 540
rect 1780 520 2280 540
rect 2320 520 2820 540
rect -1720 300 -1220 320
rect -1690 270 -1650 300
rect -1590 270 -1550 300
rect -1490 270 -1450 300
rect -1390 270 -1350 300
rect -1290 270 -1250 300
rect -1720 250 -1220 270
rect -1180 300 -680 320
rect -1150 270 -1110 300
rect -1050 270 -1010 300
rect -950 270 -910 300
rect -850 270 -810 300
rect -750 270 -710 300
rect -1180 250 -680 270
rect -540 300 -40 320
rect -510 270 -470 300
rect -410 270 -370 300
rect -310 270 -270 300
rect -210 270 -170 300
rect -110 270 -70 300
rect -540 250 -40 270
rect 0 300 500 320
rect 30 270 70 300
rect 130 270 170 300
rect 230 270 270 300
rect 330 270 370 300
rect 430 270 470 300
rect 0 250 500 270
rect 600 300 1100 320
rect 630 270 670 300
rect 730 270 770 300
rect 830 270 870 300
rect 930 270 970 300
rect 1030 270 1070 300
rect 600 250 1100 270
rect 1140 300 1640 320
rect 1170 270 1210 300
rect 1270 270 1310 300
rect 1370 270 1410 300
rect 1470 270 1510 300
rect 1570 270 1610 300
rect 1140 250 1640 270
rect 1780 300 2280 320
rect 1810 270 1850 300
rect 1910 270 1950 300
rect 2010 270 2050 300
rect 2110 270 2150 300
rect 2210 270 2250 300
rect 1780 250 2280 270
rect 2320 300 2820 320
rect 2350 270 2390 300
rect 2450 270 2490 300
rect 2550 270 2590 300
rect 2650 270 2690 300
rect 2750 270 2790 300
rect 2320 250 2820 270
rect -1720 30 -1220 50
rect -1180 30 -680 50
rect -540 30 -40 50
rect -1260 20 -1220 30
rect -1260 0 -1250 20
rect -1230 0 -1220 20
rect -1260 -10 -1220 0
rect -720 20 -680 30
rect -720 0 -710 20
rect -690 0 -680 20
rect -80 10 -70 30
rect -50 10 -40 30
rect 0 30 500 50
rect 0 10 470 30
rect 490 10 500 30
rect -80 0 -40 10
rect 460 0 500 10
rect 600 30 1100 50
rect 600 10 610 30
rect 630 10 1100 30
rect 1140 30 1640 50
rect 1780 30 2280 50
rect 2320 30 2820 50
rect 1140 10 1150 30
rect 1170 10 1180 30
rect 600 0 640 10
rect 1140 0 1180 10
rect 1780 20 1820 30
rect 1780 0 1790 20
rect 1810 0 1820 20
rect -720 -10 -680 0
rect 1780 -10 1820 0
rect 2320 20 2360 30
rect 2320 0 2330 20
rect 2350 0 2360 20
rect 2320 -10 2360 0
<< polycont >>
rect -1250 1090 -1230 1110
rect -170 1090 -150 1110
rect 1250 1090 1270 1110
rect 2330 1090 2350 1110
rect 540 970 560 990
rect -1250 0 -1230 20
rect -710 0 -690 20
rect -70 10 -50 30
rect 470 10 490 30
rect 610 10 630 30
rect 1150 10 1170 30
rect 1790 0 1810 20
rect 2330 0 2350 20
<< locali >>
rect -1260 1110 -1180 1120
rect -1260 1090 -1250 1110
rect -1230 1090 -1180 1110
rect -1260 1080 -1180 1090
rect -180 1110 1280 1120
rect -180 1090 -170 1110
rect -150 1090 1250 1110
rect 1270 1090 1280 1110
rect -180 1080 1280 1090
rect 2280 1110 2360 1120
rect 2280 1090 2330 1110
rect 2350 1090 2360 1110
rect 2280 1080 2360 1090
rect -1760 970 -1720 1060
rect -1760 950 -1750 970
rect -1730 950 -1720 970
rect -1760 860 -1720 950
rect -1790 840 -1720 860
rect -1790 810 -1780 840
rect -1760 810 -1720 840
rect -1790 790 -1720 810
rect -1760 700 -1720 790
rect -1760 680 -1750 700
rect -1730 680 -1720 700
rect -1760 580 -1720 680
rect -1220 970 -1180 1080
rect -1220 950 -1210 970
rect -1190 950 -1180 970
rect -1220 700 -1180 950
rect -1220 680 -1210 700
rect -1190 680 -1180 700
rect -1220 580 -1180 680
rect -140 1020 1240 1060
rect -140 970 -100 1020
rect 530 990 570 1000
rect 530 980 540 990
rect -140 950 -130 970
rect -110 950 -100 970
rect -140 700 -100 950
rect -140 680 -130 700
rect -110 680 -100 700
rect -140 670 -100 680
rect 400 970 540 980
rect 560 980 570 990
rect 560 970 700 980
rect 400 950 410 970
rect 430 950 670 970
rect 690 950 700 970
rect 400 940 700 950
rect 400 860 440 940
rect 660 860 700 940
rect 400 840 470 860
rect 400 810 440 840
rect 460 810 470 840
rect 400 790 470 810
rect 630 840 700 860
rect 630 810 640 840
rect 660 810 700 840
rect 630 790 700 810
rect 400 700 440 790
rect 400 680 410 700
rect 430 680 440 700
rect 400 580 440 680
rect 660 700 700 790
rect 660 680 670 700
rect 690 680 700 700
rect 660 580 700 680
rect 1200 970 1240 1020
rect 1200 950 1210 970
rect 1230 950 1240 970
rect 1200 700 1240 950
rect 1200 680 1210 700
rect 1230 680 1240 700
rect 1200 670 1240 680
rect 2280 970 2320 1080
rect 2280 950 2290 970
rect 2310 950 2320 970
rect 2280 700 2320 950
rect 2280 680 2290 700
rect 2310 680 2320 700
rect 2280 580 2320 680
rect 2820 970 2860 1060
rect 2820 950 2830 970
rect 2850 950 2860 970
rect 2820 860 2860 950
rect 2820 840 2890 860
rect 2820 810 2860 840
rect 2880 810 2890 840
rect 2820 790 2890 810
rect 2820 700 2860 790
rect 2820 680 2830 700
rect 2850 680 2860 700
rect 2820 580 2860 680
rect -1760 570 -140 580
rect -100 570 1200 580
rect 1240 570 2860 580
rect -1760 530 2860 570
rect -1760 430 -1720 530
rect -1760 410 -1750 430
rect -1730 410 -1720 430
rect -1760 320 -1720 410
rect -1790 300 -1720 320
rect -1790 270 -1780 300
rect -1760 270 -1720 300
rect -1790 250 -1720 270
rect -1760 160 -1720 250
rect -1760 140 -1750 160
rect -1730 140 -1720 160
rect -1760 50 -1720 140
rect -1220 430 -1180 530
rect -80 470 1180 510
rect -1220 410 -1210 430
rect -1190 410 -1180 430
rect -1220 160 -1180 410
rect -1220 140 -1210 160
rect -1190 140 -1180 160
rect -1220 30 -1180 140
rect -680 430 -540 440
rect -680 410 -670 430
rect -650 410 -570 430
rect -550 410 -540 430
rect -680 400 -540 410
rect -680 170 -640 400
rect -580 170 -540 400
rect -680 160 -540 170
rect -680 140 -670 160
rect -650 140 -570 160
rect -550 140 -540 160
rect -680 130 -540 140
rect -680 30 -640 130
rect -1260 20 -1180 30
rect -1260 0 -1250 20
rect -1230 0 -1180 20
rect -1260 -10 -1180 0
rect -720 20 -640 30
rect -720 0 -710 20
rect -690 0 -640 20
rect -80 30 -40 470
rect -80 10 -70 30
rect -50 10 -40 30
rect -80 0 -40 10
rect 460 410 640 450
rect 460 30 500 410
rect 460 10 470 30
rect 490 10 500 30
rect 460 0 500 10
rect 530 380 570 390
rect 530 360 540 380
rect 560 360 570 380
rect 530 300 570 360
rect 530 270 540 300
rect 560 270 570 300
rect 530 160 570 270
rect 530 140 540 160
rect 560 140 570 160
rect 530 0 570 140
rect 600 30 640 410
rect 600 10 610 30
rect 630 10 640 30
rect 600 0 640 10
rect 1140 30 1180 470
rect 1640 430 1780 440
rect 1640 410 1650 430
rect 1670 410 1750 430
rect 1770 410 1780 430
rect 1640 400 1780 410
rect 1640 170 1680 400
rect 1740 170 1780 400
rect 1640 160 1780 170
rect 1640 140 1650 160
rect 1670 140 1750 160
rect 1770 140 1780 160
rect 1640 130 1780 140
rect 1140 10 1150 30
rect 1170 10 1180 30
rect 1140 0 1180 10
rect 1740 30 1780 130
rect 2280 430 2320 530
rect 2280 410 2290 430
rect 2310 410 2320 430
rect 2280 160 2320 410
rect 2280 140 2290 160
rect 2310 140 2320 160
rect 2280 30 2320 140
rect 2820 430 2860 530
rect 2820 410 2830 430
rect 2850 410 2860 430
rect 2820 320 2860 410
rect 2820 300 2890 320
rect 2820 270 2860 300
rect 2880 270 2890 300
rect 2820 250 2890 270
rect 2820 160 2860 250
rect 2820 140 2830 160
rect 2850 140 2860 160
rect 2820 50 2860 140
rect 1740 20 1820 30
rect 1740 0 1790 20
rect 1810 0 1820 20
rect -720 -10 -640 0
rect 1740 -10 1820 0
rect 2280 20 2360 30
rect 2280 0 2330 20
rect 2350 0 2360 20
rect 2280 -10 2360 0
<< labels >>
rlabel locali -1760 550 -1760 550 7 VP
port 0 w
rlabel locali 550 0 550 0 5 VN
port 1 s
rlabel locali 480 0 480 0 5 Vdsg
port 2 s
rlabel locali -60 0 -60 0 5 Vcn
port 3 s
rlabel locali -180 1100 -180 1100 7 Vcp
port 4 w
rlabel locali -140 1040 -140 1040 7 Vout
port 5 w
<< end >>
