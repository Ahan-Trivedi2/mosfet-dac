magic
tech sky130A
timestamp 1762030467
<< error_p >>
rect 1700 1030 1718 1048
rect 1682 1010 1718 1030
rect 1700 992 1718 1010
<< nwell >>
rect -310 -90 1700 2310
<< nmos >>
rect -160 2360 -60 2460
rect -20 2360 80 2460
rect 120 2360 220 2460
rect 260 2360 360 2460
rect 400 2360 500 2460
rect 540 2360 640 2460
rect 680 2360 780 2460
rect 820 2360 920 2460
rect 960 2360 1060 2460
rect 1100 2360 1200 2460
rect 1240 2360 1340 2460
<< pmos >>
rect 0 2150 100 2250
rect 170 2150 270 2250
rect 340 2150 440 2250
rect 510 2150 610 2250
rect 680 2150 780 2250
rect 850 2150 950 2250
rect 1020 2150 1120 2250
rect 1190 2150 1290 2250
rect 1360 2150 1460 2250
rect 1530 2150 1630 2250
rect -280 1580 -80 2080
rect -280 1040 -80 1540
rect 0 1040 100 2040
rect 170 1040 270 2040
rect 340 1040 440 2040
rect 510 1040 610 2040
rect 680 1040 780 2040
rect 850 1040 950 2040
rect 1020 1040 1120 2040
rect 1190 1040 1290 2040
rect 1360 1040 1460 2040
rect 1530 1040 1630 2040
rect 0 0 100 1000
rect 170 0 270 1000
rect 340 0 440 1000
rect 510 0 610 1000
rect 680 0 780 1000
rect 850 0 950 1000
rect 1020 0 1120 1000
rect 1190 0 1290 1000
rect 1360 0 1460 1000
rect 1530 0 1630 1000
<< ndiff >>
rect 1550 2510 1700 2520
rect 1550 2490 1560 2510
rect 1580 2490 1700 2510
rect 1550 2480 1700 2490
rect -200 2430 -160 2460
rect -200 2390 -190 2430
rect -170 2390 -160 2430
rect -200 2370 -160 2390
rect -240 2360 -160 2370
rect -60 2430 -20 2460
rect -60 2390 -50 2430
rect -30 2390 -20 2430
rect -60 2360 -20 2390
rect 80 2430 120 2460
rect 80 2390 90 2430
rect 110 2390 120 2430
rect 80 2360 120 2390
rect 220 2430 260 2460
rect 220 2390 230 2430
rect 250 2390 260 2430
rect 220 2360 260 2390
rect 360 2430 400 2460
rect 360 2390 370 2430
rect 390 2390 400 2430
rect 360 2360 400 2390
rect 500 2430 540 2460
rect 500 2390 510 2430
rect 530 2390 540 2430
rect 500 2360 540 2390
rect 640 2430 680 2460
rect 640 2390 650 2430
rect 670 2390 680 2430
rect 640 2360 680 2390
rect 780 2430 820 2460
rect 780 2390 790 2430
rect 810 2390 820 2430
rect 780 2360 820 2390
rect 920 2430 960 2460
rect 920 2390 930 2430
rect 950 2390 960 2430
rect 920 2360 960 2390
rect 1060 2430 1100 2460
rect 1060 2390 1070 2430
rect 1090 2390 1100 2430
rect 1060 2360 1100 2390
rect 1200 2430 1240 2460
rect 1200 2390 1210 2430
rect 1230 2390 1240 2430
rect 1200 2360 1240 2390
rect 1340 2430 1380 2460
rect 1340 2390 1350 2430
rect 1370 2390 1380 2430
rect 1480 2440 1700 2450
rect 1480 2420 1490 2440
rect 1510 2420 1700 2440
rect 1480 2410 1520 2420
rect 1340 2360 1380 2390
rect 1550 2380 1700 2390
rect 1550 2360 1560 2380
rect 1580 2360 1700 2380
rect 1550 2350 1590 2360
<< pdiff >>
rect 0 2280 100 2290
rect 0 2260 30 2280
rect 70 2260 100 2280
rect 0 2250 100 2260
rect 170 2280 270 2290
rect 170 2260 200 2280
rect 240 2260 270 2280
rect 170 2250 270 2260
rect 340 2280 440 2290
rect 340 2260 370 2280
rect 410 2260 440 2280
rect 340 2250 440 2260
rect 510 2280 610 2290
rect 510 2260 540 2280
rect 580 2260 610 2280
rect 510 2250 610 2260
rect 680 2280 780 2290
rect 680 2260 710 2280
rect 750 2260 780 2280
rect 680 2250 780 2260
rect 850 2280 950 2290
rect 850 2260 880 2280
rect 920 2260 950 2280
rect 850 2250 950 2260
rect 1020 2280 1120 2290
rect 1020 2260 1050 2280
rect 1090 2260 1120 2280
rect 1020 2250 1120 2260
rect 1190 2280 1290 2290
rect 1190 2260 1220 2280
rect 1260 2260 1290 2280
rect 1190 2250 1290 2260
rect 1360 2280 1460 2290
rect 1360 2260 1390 2280
rect 1430 2260 1460 2280
rect 1360 2250 1460 2260
rect 1530 2280 1630 2290
rect 1530 2260 1560 2280
rect 1600 2260 1630 2280
rect 1530 2250 1630 2260
rect -280 2110 -80 2120
rect -280 2090 -200 2110
rect -160 2090 -80 2110
rect -280 2080 -80 2090
rect 0 2120 100 2150
rect 0 2070 100 2080
rect 0 2050 30 2070
rect 70 2050 100 2070
rect 0 2040 100 2050
rect 170 2120 270 2150
rect 170 2070 270 2080
rect 170 2050 200 2070
rect 240 2050 270 2070
rect 170 2040 270 2050
rect 340 2120 440 2150
rect 340 2070 440 2080
rect 340 2050 370 2070
rect 410 2050 440 2070
rect 340 2040 440 2050
rect 510 2120 610 2150
rect 510 2070 610 2080
rect 510 2050 540 2070
rect 580 2050 610 2070
rect 510 2040 610 2050
rect 680 2120 780 2150
rect 680 2070 780 2080
rect 680 2050 710 2070
rect 750 2050 780 2070
rect 680 2040 780 2050
rect 850 2120 950 2150
rect 850 2070 950 2080
rect 850 2050 880 2070
rect 920 2050 950 2070
rect 850 2040 950 2050
rect 1020 2120 1120 2150
rect 1020 2070 1120 2080
rect 1020 2050 1050 2070
rect 1090 2050 1120 2070
rect 1020 2040 1120 2050
rect 1190 2120 1290 2150
rect 1190 2070 1290 2080
rect 1190 2050 1220 2070
rect 1260 2050 1290 2070
rect 1190 2040 1290 2050
rect 1360 2120 1460 2150
rect 1360 2070 1460 2080
rect 1360 2050 1390 2070
rect 1430 2050 1460 2070
rect 1360 2040 1460 2050
rect 1530 2120 1630 2150
rect 1530 2070 1630 2080
rect 1530 2050 1560 2070
rect 1600 2050 1630 2070
rect 1530 2040 1630 2050
rect -280 1570 -80 1580
rect -280 1550 -200 1570
rect -160 1550 -80 1570
rect -280 1540 -80 1550
rect -280 1030 -80 1040
rect 0 1030 100 1040
rect 170 1030 270 1040
rect 340 1030 440 1040
rect 510 1030 610 1040
rect 680 1030 780 1040
rect 850 1030 950 1040
rect 1020 1030 1120 1040
rect 1190 1030 1290 1040
rect 1360 1030 1460 1040
rect 1530 1030 1630 1040
rect -280 1010 -200 1030
rect -160 1010 30 1030
rect 70 1010 200 1030
rect 240 1010 370 1030
rect 410 1010 540 1030
rect 580 1010 710 1030
rect 750 1010 880 1030
rect 920 1010 1050 1030
rect 1090 1010 1220 1030
rect 1260 1010 1390 1030
rect 1430 1010 1560 1030
rect 1600 1010 1700 1030
rect -280 1000 -80 1010
rect 0 1000 100 1010
rect 170 1000 270 1010
rect 340 1000 440 1010
rect 510 1000 610 1010
rect 680 1000 780 1010
rect 850 1000 950 1010
rect 1020 1000 1120 1010
rect 1190 1000 1290 1010
rect 1360 1000 1460 1010
rect 1530 1000 1630 1010
rect 0 -10 100 0
rect 0 -30 30 -10
rect 70 -30 100 -10
rect 0 -40 100 -30
rect 170 -10 270 0
rect 170 -30 200 -10
rect 240 -30 270 -10
rect 170 -40 270 -30
rect 340 -10 440 0
rect 340 -30 370 -10
rect 410 -30 440 -10
rect 340 -40 440 -30
rect 510 -10 610 0
rect 510 -30 540 -10
rect 580 -30 610 -10
rect 510 -40 610 -30
rect 680 -10 780 0
rect 680 -30 710 -10
rect 750 -30 780 -10
rect 680 -40 780 -30
rect 850 -10 950 0
rect 850 -30 880 -10
rect 920 -30 950 -10
rect 850 -40 950 -30
rect 1020 -10 1120 0
rect 1020 -30 1050 -10
rect 1090 -30 1120 -10
rect 1020 -40 1120 -30
rect 1190 -10 1290 0
rect 1190 -30 1220 -10
rect 1260 -30 1290 -10
rect 1190 -40 1290 -30
rect 1360 -10 1460 0
rect 1360 -30 1390 -10
rect 1430 -30 1460 -10
rect 1360 -40 1460 -30
rect 1530 -10 1630 0
rect 1530 -30 1560 -10
rect 1600 -30 1630 -10
rect 1530 -40 1630 -30
<< ndiffc >>
rect 1560 2490 1580 2510
rect -190 2390 -170 2430
rect -50 2390 -30 2430
rect 90 2390 110 2430
rect 230 2390 250 2430
rect 370 2390 390 2430
rect 510 2390 530 2430
rect 650 2390 670 2430
rect 790 2390 810 2430
rect 930 2390 950 2430
rect 1070 2390 1090 2430
rect 1210 2390 1230 2430
rect 1350 2390 1370 2430
rect 1490 2420 1510 2440
rect 1560 2360 1580 2380
<< pdiffc >>
rect 30 2260 70 2280
rect 200 2260 240 2280
rect 370 2260 410 2280
rect 540 2260 580 2280
rect 710 2260 750 2280
rect 880 2260 920 2280
rect 1050 2260 1090 2280
rect 1220 2260 1260 2280
rect 1390 2260 1430 2280
rect 1560 2260 1600 2280
rect -200 2090 -160 2110
rect 30 2050 70 2070
rect 200 2050 240 2070
rect 370 2050 410 2070
rect 540 2050 580 2070
rect 710 2050 750 2070
rect 880 2050 920 2070
rect 1050 2050 1090 2070
rect 1220 2050 1260 2070
rect 1390 2050 1430 2070
rect 1560 2050 1600 2070
rect -200 1550 -160 1570
rect -200 1010 -160 1030
rect 30 1010 70 1030
rect 200 1010 240 1030
rect 370 1010 410 1030
rect 540 1010 580 1030
rect 710 1010 750 1030
rect 880 1010 920 1030
rect 1050 1010 1090 1030
rect 1220 1010 1260 1030
rect 1390 1010 1430 1030
rect 1560 1010 1600 1030
rect 30 -30 70 -10
rect 200 -30 240 -10
rect 370 -30 410 -10
rect 540 -30 580 -10
rect 710 -30 750 -10
rect 880 -30 920 -10
rect 1050 -30 1090 -10
rect 1220 -30 1260 -10
rect 1390 -30 1430 -10
rect 1560 -30 1600 -10
<< psubdiff >>
rect 1400 2500 1460 2520
rect 1400 2480 1420 2500
rect 1440 2480 1460 2500
rect 1410 2470 1450 2480
rect -240 2430 -200 2460
rect -240 2390 -230 2430
rect -210 2390 -200 2430
rect -240 2370 -200 2390
<< nsubdiff >>
rect 0 2110 100 2120
rect 0 2090 30 2110
rect 70 2090 100 2110
rect 0 2080 100 2090
rect 170 2110 270 2120
rect 170 2090 200 2110
rect 240 2090 270 2110
rect 170 2080 270 2090
rect 340 2110 440 2120
rect 340 2090 370 2110
rect 410 2090 440 2110
rect 340 2080 440 2090
rect 510 2110 610 2120
rect 510 2090 540 2110
rect 580 2090 610 2110
rect 510 2080 610 2090
rect 680 2110 780 2120
rect 680 2090 710 2110
rect 750 2090 780 2110
rect 680 2080 780 2090
rect 850 2110 950 2120
rect 850 2090 880 2110
rect 920 2090 950 2110
rect 850 2080 950 2090
rect 1020 2110 1120 2120
rect 1020 2090 1050 2110
rect 1090 2090 1120 2110
rect 1020 2080 1120 2090
rect 1190 2110 1290 2120
rect 1190 2090 1220 2110
rect 1260 2090 1290 2110
rect 1190 2080 1290 2090
rect 1360 2110 1460 2120
rect 1360 2090 1390 2110
rect 1430 2090 1460 2110
rect 1360 2080 1460 2090
rect 1530 2110 1630 2120
rect 1530 2090 1560 2110
rect 1600 2090 1630 2110
rect 1530 2080 1630 2090
rect 0 -50 100 -40
rect 0 -70 30 -50
rect 70 -70 100 -50
rect 170 -50 270 -40
rect 170 -70 200 -50
rect 240 -70 270 -50
rect 340 -50 440 -40
rect 340 -70 370 -50
rect 410 -70 440 -50
rect 510 -50 610 -40
rect 510 -70 540 -50
rect 580 -70 610 -50
rect 680 -50 780 -40
rect 680 -70 710 -50
rect 750 -70 780 -50
rect 850 -50 950 -40
rect 850 -70 880 -50
rect 920 -70 950 -50
rect 1020 -50 1120 -40
rect 1020 -70 1050 -50
rect 1090 -70 1120 -50
rect 1190 -50 1290 -40
rect 1190 -70 1220 -50
rect 1260 -70 1290 -50
rect 1360 -50 1460 -40
rect 1360 -70 1390 -50
rect 1430 -70 1460 -50
rect 1530 -50 1630 -40
rect 1530 -70 1560 -50
rect 1600 -70 1630 -50
<< psubdiffcont >>
rect 1420 2480 1440 2500
rect -230 2390 -210 2430
<< nsubdiffcont >>
rect 30 2090 70 2110
rect 200 2090 240 2110
rect 370 2090 410 2110
rect 540 2090 580 2110
rect 710 2090 750 2110
rect 880 2090 920 2110
rect 1050 2090 1090 2110
rect 1220 2090 1260 2110
rect 1390 2090 1430 2110
rect 1560 2090 1600 2110
rect 30 -70 70 -50
rect 200 -70 240 -50
rect 370 -70 410 -50
rect 540 -70 580 -50
rect 710 -70 750 -50
rect 880 -70 920 -50
rect 1050 -70 1090 -50
rect 1220 -70 1260 -50
rect 1390 -70 1430 -50
rect 1560 -70 1600 -50
<< poly >>
rect -160 2460 -60 2480
rect -20 2460 80 2480
rect 120 2460 220 2480
rect 260 2460 360 2480
rect 400 2460 500 2480
rect 540 2460 640 2480
rect 680 2460 780 2480
rect 820 2460 920 2480
rect 960 2460 1060 2480
rect 1100 2460 1200 2480
rect 1240 2460 1340 2480
rect -160 2350 -60 2360
rect -200 2340 -60 2350
rect -20 2350 80 2360
rect 120 2350 220 2360
rect -20 2340 220 2350
rect 260 2350 360 2360
rect 400 2350 500 2360
rect 260 2340 500 2350
rect 540 2350 640 2360
rect 680 2350 780 2360
rect 540 2340 780 2350
rect 820 2350 920 2360
rect 960 2350 1060 2360
rect 820 2340 1060 2350
rect 1100 2350 1200 2360
rect 1240 2350 1340 2360
rect 1100 2340 1340 2350
rect 1610 2340 1660 2350
rect -200 2320 -190 2340
rect -170 2330 -140 2340
rect 60 2330 90 2340
rect -170 2320 -160 2330
rect -200 2310 -160 2320
rect 80 2320 90 2330
rect 110 2330 140 2340
rect 340 2330 370 2340
rect 110 2320 120 2330
rect 80 2310 120 2320
rect 360 2320 370 2330
rect 390 2330 420 2340
rect 620 2330 650 2340
rect 390 2320 400 2330
rect 360 2310 400 2320
rect 640 2320 650 2330
rect 670 2330 700 2340
rect 900 2330 930 2340
rect 670 2320 680 2330
rect 640 2310 680 2320
rect 920 2320 930 2330
rect 950 2330 980 2340
rect 1180 2330 1210 2340
rect 950 2320 960 2330
rect 920 2310 960 2320
rect 1200 2320 1210 2330
rect 1230 2330 1260 2340
rect 1230 2320 1240 2330
rect 1200 2310 1240 2320
rect 1610 2320 1620 2340
rect 1640 2320 1660 2340
rect 1610 2310 1660 2320
rect 1640 2250 1660 2310
rect -90 2170 -50 2180
rect -90 2150 -80 2170
rect -60 2150 -50 2170
rect -20 2150 0 2250
rect 100 2210 120 2250
rect 150 2210 170 2250
rect 100 2190 170 2210
rect 100 2150 120 2190
rect 150 2150 170 2190
rect 270 2210 290 2250
rect 320 2210 340 2250
rect 270 2190 340 2210
rect 270 2150 290 2190
rect 320 2150 340 2190
rect 440 2210 460 2250
rect 490 2210 510 2250
rect 440 2190 510 2210
rect 440 2150 460 2190
rect 490 2150 510 2190
rect 610 2210 630 2250
rect 660 2210 680 2250
rect 610 2190 680 2210
rect 610 2150 630 2190
rect 660 2150 680 2190
rect 780 2210 800 2250
rect 830 2210 850 2250
rect 780 2190 850 2210
rect 780 2150 800 2190
rect 830 2150 850 2190
rect 950 2210 970 2250
rect 1000 2210 1020 2250
rect 950 2190 1020 2210
rect 950 2150 970 2190
rect 1000 2150 1020 2190
rect 1120 2210 1140 2250
rect 1170 2210 1190 2250
rect 1120 2190 1190 2210
rect 1120 2150 1140 2190
rect 1170 2150 1190 2190
rect 1290 2210 1310 2250
rect 1340 2210 1360 2250
rect 1290 2190 1360 2210
rect 1290 2150 1310 2190
rect 1340 2150 1360 2190
rect 1460 2210 1480 2250
rect 1510 2210 1530 2250
rect 1460 2190 1530 2210
rect 1460 2150 1480 2190
rect 1510 2150 1530 2190
rect 1630 2210 1660 2250
rect 1630 2190 1700 2210
rect 1630 2150 1650 2190
rect -90 2140 -50 2150
rect -70 2080 -50 2140
rect -300 1580 -280 2080
rect -80 2060 -50 2080
rect -80 1580 -60 2060
rect -300 1060 -280 1540
rect -310 1040 -280 1060
rect -80 1040 -60 1540
rect -20 1040 0 2040
rect 100 1550 120 2040
rect 150 1550 170 2040
rect 100 1530 170 1550
rect 100 1040 120 1530
rect 150 1040 170 1530
rect 270 1550 290 2040
rect 320 1550 340 2040
rect 270 1530 340 1550
rect 270 1040 290 1530
rect 320 1040 340 1530
rect 440 1550 460 2040
rect 490 1550 510 2040
rect 440 1530 510 1550
rect 440 1040 460 1530
rect 490 1040 510 1530
rect 610 1550 630 2040
rect 660 1550 680 2040
rect 610 1530 680 1550
rect 610 1040 630 1530
rect 660 1040 680 1530
rect 780 1550 800 2040
rect 830 1550 850 2040
rect 780 1530 850 1550
rect 780 1040 800 1530
rect 830 1040 850 1530
rect 950 1550 970 2040
rect 1000 1550 1020 2040
rect 950 1530 1020 1550
rect 950 1040 970 1530
rect 1000 1040 1020 1530
rect 1120 1550 1140 2040
rect 1170 1550 1190 2040
rect 1120 1530 1190 1550
rect 1120 1040 1140 1530
rect 1170 1040 1190 1530
rect 1290 1550 1310 2040
rect 1340 1550 1360 2040
rect 1290 1530 1360 1550
rect 1290 1040 1310 1530
rect 1340 1040 1360 1530
rect 1460 1550 1480 2040
rect 1510 1550 1530 2040
rect 1460 1530 1530 1550
rect 1460 1040 1480 1530
rect 1510 1040 1530 1530
rect 1630 1550 1650 2040
rect 1630 1530 1700 1550
rect 1630 1040 1650 1530
rect -310 980 -290 1040
rect -310 970 -270 980
rect -310 950 -300 970
rect -280 950 -270 970
rect -310 940 -270 950
rect -20 0 0 1000
rect 100 510 120 1000
rect 150 510 170 1000
rect 100 490 170 510
rect 100 0 120 490
rect 150 0 170 490
rect 270 510 290 1000
rect 320 510 340 1000
rect 270 490 340 510
rect 270 0 290 490
rect 320 0 340 490
rect 440 510 460 1000
rect 490 510 510 1000
rect 440 490 510 510
rect 440 0 460 490
rect 490 0 510 490
rect 610 510 630 1000
rect 660 510 680 1000
rect 610 490 680 510
rect 610 0 630 490
rect 660 0 680 490
rect 780 510 800 1000
rect 830 510 850 1000
rect 780 490 850 510
rect 780 0 800 490
rect 830 0 850 490
rect 950 510 970 1000
rect 1000 510 1020 1000
rect 950 490 1020 510
rect 950 0 970 490
rect 1000 0 1020 490
rect 1120 510 1140 1000
rect 1170 510 1190 1000
rect 1120 490 1190 510
rect 1120 0 1140 490
rect 1170 0 1190 490
rect 1290 510 1310 1000
rect 1340 510 1360 1000
rect 1290 490 1360 510
rect 1290 0 1310 490
rect 1340 0 1360 490
rect 1460 510 1480 1000
rect 1510 510 1530 1000
rect 1460 490 1530 510
rect 1460 0 1480 490
rect 1510 0 1530 490
rect 1630 510 1650 1000
rect 1630 490 1700 510
rect 1630 0 1650 490
<< polycont >>
rect -190 2320 -170 2340
rect 90 2320 110 2340
rect 370 2320 390 2340
rect 650 2320 670 2340
rect 930 2320 950 2340
rect 1210 2320 1230 2340
rect 1620 2320 1640 2340
rect -80 2150 -60 2170
rect -300 950 -280 970
<< locali >>
rect -190 2510 1590 2520
rect -190 2500 1560 2510
rect -190 2440 -170 2500
rect 1410 2480 1420 2500
rect 1440 2480 1450 2500
rect 1550 2490 1560 2500
rect 1580 2490 1590 2510
rect 1550 2480 1590 2490
rect -50 2460 1370 2480
rect 1410 2470 1450 2480
rect -50 2440 -30 2460
rect 230 2440 250 2460
rect 510 2440 530 2460
rect 790 2440 810 2460
rect 1070 2440 1090 2460
rect 1350 2440 1370 2460
rect 1480 2440 1520 2450
rect -240 2430 -160 2440
rect -240 2390 -230 2430
rect -210 2390 -190 2430
rect -170 2390 -160 2430
rect -240 2380 -160 2390
rect -60 2430 -20 2440
rect -60 2390 -50 2430
rect -30 2390 -20 2430
rect -60 2380 -20 2390
rect 80 2430 120 2440
rect 80 2390 90 2430
rect 110 2390 120 2430
rect 80 2380 120 2390
rect 220 2430 260 2440
rect 220 2390 230 2430
rect 250 2390 260 2430
rect 220 2380 260 2390
rect 360 2430 400 2440
rect 360 2390 370 2430
rect 390 2390 400 2430
rect 360 2380 400 2390
rect 500 2430 540 2440
rect 500 2390 510 2430
rect 530 2390 540 2430
rect 500 2380 540 2390
rect 640 2430 680 2440
rect 640 2390 650 2430
rect 670 2390 680 2430
rect 640 2380 680 2390
rect 780 2430 820 2440
rect 780 2390 790 2430
rect 810 2390 820 2430
rect 780 2380 820 2390
rect 920 2430 960 2440
rect 920 2390 930 2430
rect 950 2390 960 2430
rect 920 2380 960 2390
rect 1060 2430 1100 2440
rect 1060 2390 1070 2430
rect 1090 2390 1100 2430
rect 1060 2380 1100 2390
rect 1200 2430 1240 2440
rect 1200 2390 1210 2430
rect 1230 2390 1240 2430
rect 1200 2380 1240 2390
rect 1340 2430 1490 2440
rect 1340 2390 1350 2430
rect 1370 2420 1490 2430
rect 1510 2420 1520 2440
rect 1370 2390 1380 2420
rect 1480 2410 1520 2420
rect 1340 2380 1380 2390
rect 1550 2380 1590 2390
rect -190 2350 -170 2380
rect -200 2340 -160 2350
rect -200 2320 -190 2340
rect -170 2320 -160 2340
rect -50 2320 -30 2380
rect 90 2350 110 2380
rect 370 2350 390 2380
rect 650 2350 670 2380
rect 930 2350 950 2380
rect 1210 2350 1230 2380
rect 1550 2360 1560 2380
rect 1580 2360 1590 2380
rect 1550 2350 1590 2360
rect 1620 2350 1640 2520
rect -200 2310 -160 2320
rect -190 2120 -170 2310
rect -130 2300 -30 2320
rect 80 2340 120 2350
rect 360 2340 400 2350
rect 640 2340 680 2350
rect 920 2340 960 2350
rect 1200 2340 1240 2350
rect 1550 2340 1570 2350
rect 80 2320 90 2340
rect 110 2320 370 2340
rect 390 2320 650 2340
rect 670 2320 930 2340
rect 950 2320 1210 2340
rect 1230 2320 1570 2340
rect 1610 2340 1650 2350
rect 1610 2320 1620 2340
rect 1640 2320 1650 2340
rect 80 2310 120 2320
rect 360 2310 400 2320
rect 640 2310 680 2320
rect 920 2310 960 2320
rect 1200 2310 1240 2320
rect 1610 2310 1650 2320
rect -210 2110 -150 2120
rect -210 2090 -200 2110
rect -160 2090 -150 2110
rect -210 2080 -150 2090
rect -210 1570 -150 1580
rect -130 1570 -110 2300
rect 20 2280 80 2290
rect 190 2280 250 2290
rect 360 2280 420 2290
rect 530 2280 590 2290
rect 700 2280 760 2290
rect 870 2280 930 2290
rect 1040 2280 1100 2290
rect 1210 2280 1270 2290
rect 1380 2280 1440 2290
rect 1550 2280 1610 2290
rect -80 2260 30 2280
rect 70 2260 200 2280
rect 240 2260 370 2280
rect 410 2260 540 2280
rect 580 2260 710 2280
rect 750 2260 880 2280
rect 920 2260 1050 2280
rect 1090 2260 1220 2280
rect 1260 2260 1390 2280
rect 1430 2260 1560 2280
rect 1600 2260 1610 2280
rect -80 2180 -60 2260
rect 20 2250 80 2260
rect 190 2250 250 2260
rect 360 2250 420 2260
rect 530 2250 590 2260
rect 700 2250 760 2260
rect 870 2250 930 2260
rect 1040 2250 1100 2260
rect 1210 2250 1270 2260
rect 1380 2250 1440 2260
rect 1550 2250 1610 2260
rect -90 2170 -50 2180
rect -90 2150 -80 2170
rect -60 2150 -50 2170
rect -90 2140 -50 2150
rect 20 2110 80 2120
rect 20 2090 30 2110
rect 70 2090 80 2110
rect 190 2110 250 2120
rect 190 2090 200 2110
rect 240 2090 250 2110
rect 360 2110 420 2120
rect 360 2090 370 2110
rect 410 2090 420 2110
rect 530 2110 590 2120
rect 530 2090 540 2110
rect 580 2090 590 2110
rect 700 2110 760 2120
rect 700 2090 710 2110
rect 750 2090 760 2110
rect 870 2110 930 2120
rect 870 2090 880 2110
rect 920 2090 930 2110
rect 1040 2110 1100 2120
rect 1040 2090 1050 2110
rect 1090 2090 1100 2110
rect 1210 2110 1270 2120
rect 1210 2090 1220 2110
rect 1260 2090 1270 2110
rect 1380 2110 1440 2120
rect 1380 2090 1390 2110
rect 1430 2090 1440 2110
rect 1550 2110 1610 2120
rect 1550 2090 1560 2110
rect 1600 2090 1610 2110
rect 1680 2090 1700 2520
rect 20 2070 1700 2090
rect 20 2050 30 2070
rect 70 2050 80 2070
rect 20 2040 80 2050
rect 190 2050 200 2070
rect 240 2050 250 2070
rect 190 2040 250 2050
rect 360 2050 370 2070
rect 410 2050 420 2070
rect 360 2040 420 2050
rect 530 2050 540 2070
rect 580 2050 590 2070
rect 530 2040 590 2050
rect 700 2050 710 2070
rect 750 2050 760 2070
rect 700 2040 760 2050
rect 870 2050 880 2070
rect 920 2050 930 2070
rect 870 2040 930 2050
rect 1040 2050 1050 2070
rect 1090 2050 1100 2070
rect 1040 2040 1100 2050
rect 1210 2050 1220 2070
rect 1260 2050 1270 2070
rect 1210 2040 1270 2050
rect 1380 2050 1390 2070
rect 1430 2050 1440 2070
rect 1380 2040 1440 2050
rect 1550 2050 1560 2070
rect 1600 2050 1610 2070
rect 1550 2040 1610 2050
rect -210 1550 -200 1570
rect -160 1550 -110 1570
rect -210 1540 -150 1550
rect -210 1030 -150 1040
rect -210 1010 -200 1030
rect -160 1010 -150 1030
rect -210 1000 -150 1010
rect 20 1030 80 1040
rect 20 1010 30 1030
rect 70 1010 80 1030
rect 20 1000 80 1010
rect 190 1030 250 1040
rect 190 1010 200 1030
rect 240 1010 250 1030
rect 190 1000 250 1010
rect 360 1030 420 1040
rect 360 1010 370 1030
rect 410 1010 420 1030
rect 360 1000 420 1010
rect 530 1030 590 1040
rect 530 1010 540 1030
rect 580 1010 590 1030
rect 530 1000 590 1010
rect 700 1030 760 1040
rect 700 1010 710 1030
rect 750 1010 760 1030
rect 700 1000 760 1010
rect 870 1030 930 1040
rect 870 1010 880 1030
rect 920 1010 930 1030
rect 870 1000 930 1010
rect 1040 1030 1100 1040
rect 1040 1010 1050 1030
rect 1090 1010 1100 1030
rect 1040 1000 1100 1010
rect 1210 1030 1270 1040
rect 1210 1010 1220 1030
rect 1260 1010 1270 1030
rect 1210 1000 1270 1010
rect 1380 1030 1440 1040
rect 1380 1010 1390 1030
rect 1430 1010 1440 1030
rect 1380 1000 1440 1010
rect 1550 1030 1610 1040
rect 1550 1010 1560 1030
rect 1600 1010 1610 1030
rect 1550 1000 1610 1010
rect -310 970 -270 980
rect -190 970 -170 1000
rect -310 950 -300 970
rect -280 950 -170 970
rect -310 940 -270 950
rect 20 -10 80 0
rect 20 -30 30 -10
rect 70 -30 80 -10
rect 190 -10 250 0
rect 190 -30 200 -10
rect 240 -30 250 -10
rect 360 -10 420 0
rect 360 -30 370 -10
rect 410 -30 420 -10
rect 530 -10 590 0
rect 530 -30 540 -10
rect 580 -30 590 -10
rect 700 -10 760 0
rect 700 -30 710 -10
rect 750 -30 760 -10
rect 870 -10 930 0
rect 870 -30 880 -10
rect 920 -30 930 -10
rect 1040 -10 1100 0
rect 1040 -30 1050 -10
rect 1090 -30 1100 -10
rect 1210 -10 1270 0
rect 1210 -30 1220 -10
rect 1260 -30 1270 -10
rect 1380 -10 1440 0
rect 1380 -30 1390 -10
rect 1430 -30 1440 -10
rect 1550 -10 1610 0
rect 1550 -30 1560 -10
rect 1600 -30 1610 -10
rect 1680 -30 1700 2070
rect 20 -50 1700 -30
rect 20 -70 30 -50
rect 70 -70 80 -50
rect 190 -70 200 -50
rect 240 -70 250 -50
rect 360 -70 370 -50
rect 410 -70 420 -50
rect 530 -70 540 -50
rect 580 -70 590 -50
rect 700 -70 710 -50
rect 750 -70 760 -50
rect 870 -70 880 -50
rect 920 -70 930 -50
rect 1040 -70 1050 -50
rect 1090 -70 1100 -50
rect 1210 -70 1220 -50
rect 1260 -70 1270 -50
rect 1380 -70 1390 -50
rect 1430 -70 1440 -50
rect 1550 -70 1560 -50
rect 1600 -70 1610 -50
<< end >>
