* SPICE3 file created from ncbc.ext - technology: sky130A


* Top level circuit ncbc

X0 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X1 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X2 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X3 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X4 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X5 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X6 a_n560_3080# a_n620_1880# a_n620_1880# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X7 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X8 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X9 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X10 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X11 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X12 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X13 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X14 a_n620_1880# a_n620_1880# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X15 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X16 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X17 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X18 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X19 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X20 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X21 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X22 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X23 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X24 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X25 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X26 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X27 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X28 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X29 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X30 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X31 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X32 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X33 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X34 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X35 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X36 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X37 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X38 a_n620_1880# a_n620_1880# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X39 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X40 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X41 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X42 a_n560_3080# a_n560_4160# a_n560_4160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X43 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X44 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X45 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X46 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X47 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X48 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X49 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X50 a_n560_4160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X51 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X52 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X53 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X54 a_n560_3080# a_n600_3160# a_n560_4160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X55 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X56 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X57 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X58 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X59 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X60 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X61 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X62 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X63 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X64 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X65 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X66 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X67 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X68 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X69 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X70 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X71 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X72 a_n560_4160# a_n560_4160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X73 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X74 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X75 a_n560_3080# a_n620_1880# a_n620_1880# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X76 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X77 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X78 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X79 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X80 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X81 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X82 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X83 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X84 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X85 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X86 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X87 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X88 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X89 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X90 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X91 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X92 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X93 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X94 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X95 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X96 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X97 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X98 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X99 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X100 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X101 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X102 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X103 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X104 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X105 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X106 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X107 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X108 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X109 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X110 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X111 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X112 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X113 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X114 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X115 a_n560_4160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X116 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X117 a_n560_3080# a_n600_3160# a_n560_4160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X118 a_n560_3080# a_n560_4160# a_n560_4160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X119 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X120 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X121 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X122 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X123 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X124 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X125 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X126 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X127 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X128 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X129 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X130 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X131 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X132 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X133 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X134 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X135 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X136 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X137 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X138 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X139 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X140 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X141 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X142 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X143 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X144 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X145 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X146 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X147 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X148 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X149 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X150 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X151 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X152 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X153 a_n560_4160# a_n560_4160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X154 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X155 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X156 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X157 a_n600_3160# a_n600_3160# a_n560_3080# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X158 w_n40_1620# w_n40_1620# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X159 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X160 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X161 w_n40_1620# a_n40_2080# a_n600_3160# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X162 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X163 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X164 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X165 a_n600_3160# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X166 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X167 w_n40_1620# a_n40_2080# a_n620_1880# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X168 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X169 a_n560_3080# a_n600_3160# a_n600_3160# a_n560_4160# sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X170 a_n620_1880# w_n40_1620# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X171 a_n620_1880# a_n40_2080# w_n40_1620# w_n40_1620# sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
.end

