magic
tech sky130A
timestamp 1762047425
<< nwell >>
rect -150 -160 325 200
rect 2650 -195 3125 165
<< nmos >>
rect 415 55 915 255
rect 965 55 1465 255
rect 1515 55 2015 255
rect 2065 55 2565 255
rect 415 -365 915 -165
rect 965 -365 1465 -165
rect 1515 -365 2015 -165
rect 2065 -365 2565 -165
<< pmos >>
rect 5 80 105 180
rect 155 80 255 180
rect 2805 45 2905 145
rect 2955 45 3055 145
rect 5 -140 105 -40
rect 155 -140 255 -40
rect 2805 -175 2905 -75
rect 2955 -175 3055 -75
<< ndiff >>
rect 365 240 415 255
rect 365 70 380 240
rect 400 70 415 240
rect 365 55 415 70
rect 915 240 965 255
rect 915 70 930 240
rect 950 70 965 240
rect 915 55 965 70
rect 1465 240 1515 255
rect 1465 70 1480 240
rect 1500 70 1515 240
rect 1465 55 1515 70
rect 2015 240 2065 255
rect 2015 70 2030 240
rect 2050 70 2065 240
rect 2015 55 2065 70
rect 2565 240 2615 255
rect 2565 70 2580 240
rect 2600 70 2615 240
rect 2565 55 2615 70
rect 365 -180 415 -165
rect 365 -350 380 -180
rect 400 -350 415 -180
rect 365 -365 415 -350
rect 915 -180 965 -165
rect 915 -350 930 -180
rect 950 -350 965 -180
rect 915 -365 965 -350
rect 1465 -180 1515 -165
rect 1465 -350 1480 -180
rect 1500 -350 1515 -180
rect 1465 -365 1515 -350
rect 2015 -180 2065 -165
rect 2015 -350 2030 -180
rect 2050 -350 2065 -180
rect 2015 -365 2065 -350
rect 2565 -180 2615 -165
rect 2565 -350 2580 -180
rect 2600 -350 2615 -180
rect 2565 -365 2615 -350
<< pdiff >>
rect -45 165 5 180
rect -45 95 -30 165
rect -10 95 5 165
rect -45 80 5 95
rect 105 165 155 180
rect 105 95 120 165
rect 140 95 155 165
rect 105 80 155 95
rect 255 165 305 180
rect 255 95 270 165
rect 290 95 305 165
rect 255 80 305 95
rect 2755 130 2805 145
rect 2755 60 2770 130
rect 2790 60 2805 130
rect 2755 45 2805 60
rect 2905 130 2955 145
rect 2905 60 2920 130
rect 2940 60 2955 130
rect 2905 45 2955 60
rect 3055 130 3105 145
rect 3055 60 3070 130
rect 3090 60 3105 130
rect 3055 45 3105 60
rect -45 -55 5 -40
rect -45 -125 -30 -55
rect -10 -125 5 -55
rect -45 -140 5 -125
rect 105 -55 155 -40
rect 105 -125 120 -55
rect 140 -125 155 -55
rect 105 -140 155 -125
rect 255 -55 305 -40
rect 255 -125 270 -55
rect 290 -125 305 -55
rect 255 -140 305 -125
rect 2755 -90 2805 -75
rect 2755 -160 2770 -90
rect 2790 -160 2805 -90
rect 2755 -175 2805 -160
rect 2905 -90 2955 -75
rect 2905 -160 2920 -90
rect 2940 -160 2955 -90
rect 2905 -175 2955 -160
rect 3055 -90 3105 -75
rect 3055 -160 3070 -90
rect 3090 -160 3105 -90
rect 3055 -175 3105 -160
<< ndiffc >>
rect 380 70 400 240
rect 930 70 950 240
rect 1480 70 1500 240
rect 2030 70 2050 240
rect 2580 70 2600 240
rect 380 -350 400 -180
rect 930 -350 950 -180
rect 1480 -350 1500 -180
rect 2030 -350 2050 -180
rect 2580 -350 2600 -180
<< pdiffc >>
rect -30 95 -10 165
rect 120 95 140 165
rect 270 95 290 165
rect 2770 60 2790 130
rect 2920 60 2940 130
rect 3070 60 3090 130
rect -30 -125 -10 -55
rect 120 -125 140 -55
rect 270 -125 290 -55
rect 2770 -160 2790 -90
rect 2920 -160 2940 -90
rect 3070 -160 3090 -90
<< psubdiff >>
rect 1530 -20 1580 -5
rect 1530 -90 1545 -20
rect 1565 -90 1580 -20
rect 1530 -105 1580 -90
<< nsubdiff >>
rect -130 -55 -80 -40
rect -130 -125 -115 -55
rect -95 -125 -80 -55
rect -130 -140 -80 -125
rect 2670 -90 2720 -75
rect 2670 -160 2685 -90
rect 2705 -160 2720 -90
rect 2670 -175 2720 -160
<< psubdiffcont >>
rect 1545 -90 1565 -20
<< nsubdiffcont >>
rect -115 -125 -95 -55
rect 2685 -160 2705 -90
<< poly >>
rect 980 300 1020 310
rect 980 280 990 300
rect 1010 280 1020 300
rect 980 270 1020 280
rect 1610 300 1650 310
rect 1610 280 1620 300
rect 1640 280 1650 300
rect 1610 270 1650 280
rect 415 255 915 270
rect 965 255 1465 270
rect 1515 255 2015 270
rect 2065 255 2565 270
rect 5 180 105 195
rect 155 180 255 195
rect 5 65 105 80
rect 155 65 255 80
rect 20 55 60 65
rect 20 35 30 55
rect 50 35 60 55
rect 20 25 60 35
rect 170 55 210 65
rect 2805 145 2905 160
rect 2955 145 3055 160
rect 170 35 180 55
rect 200 35 210 55
rect 415 40 915 55
rect 965 40 1465 55
rect 1515 40 2015 55
rect 2065 40 2565 55
rect 170 25 210 35
rect 430 30 470 40
rect 430 10 440 30
rect 460 10 470 30
rect 430 0 470 10
rect 2080 30 2120 40
rect 2805 30 2905 45
rect 2955 30 3055 45
rect 2080 10 2090 30
rect 2110 10 2120 30
rect 2080 0 2120 10
rect 2820 20 2860 30
rect 2820 0 2830 20
rect 2850 0 2860 20
rect 2820 -10 2860 0
rect 2970 20 3010 30
rect 2970 0 2980 20
rect 3000 0 3010 20
rect 2970 -10 3010 0
rect 5 -40 105 -25
rect 155 -40 255 -25
rect 2805 -75 2905 -60
rect 2955 -75 3055 -60
rect 980 -120 1020 -110
rect 980 -140 990 -120
rect 1010 -140 1020 -120
rect 5 -155 105 -140
rect 155 -155 255 -140
rect 980 -150 1020 -140
rect 1610 -120 1650 -110
rect 1610 -140 1620 -120
rect 1640 -140 1650 -120
rect 1610 -150 1650 -140
rect 20 -165 60 -155
rect 20 -185 30 -165
rect 50 -185 60 -165
rect 20 -195 60 -185
rect 170 -165 210 -155
rect 415 -165 915 -150
rect 965 -165 1465 -150
rect 1515 -165 2015 -150
rect 2065 -165 2565 -150
rect 170 -185 180 -165
rect 200 -185 210 -165
rect 170 -195 210 -185
rect 2805 -190 2905 -175
rect 2955 -190 3055 -175
rect 2820 -200 2860 -190
rect 2820 -220 2830 -200
rect 2850 -220 2860 -200
rect 2820 -230 2860 -220
rect 2970 -200 3010 -190
rect 2970 -220 2980 -200
rect 3000 -220 3010 -200
rect 2970 -230 3010 -220
rect 415 -380 915 -365
rect 965 -380 1465 -365
rect 1515 -380 2015 -365
rect 2065 -380 2565 -365
rect 430 -390 470 -380
rect 430 -410 440 -390
rect 460 -410 470 -390
rect 430 -420 470 -410
rect 2080 -390 2120 -380
rect 2080 -410 2090 -390
rect 2110 -410 2120 -390
rect 2080 -420 2120 -410
<< polycont >>
rect 990 280 1010 300
rect 1620 280 1640 300
rect 30 35 50 55
rect 180 35 200 55
rect 440 10 460 30
rect 2090 10 2110 30
rect 2830 0 2850 20
rect 2980 0 3000 20
rect 990 -140 1010 -120
rect 1620 -140 1640 -120
rect 30 -185 50 -165
rect 180 -185 200 -165
rect 2830 -220 2850 -200
rect 2980 -220 3000 -200
rect 440 -410 460 -390
rect 2090 -410 2110 -390
<< locali >>
rect 120 380 2940 400
rect 120 175 140 380
rect 380 340 2595 360
rect 380 335 1010 340
rect 380 250 400 335
rect 990 310 1010 335
rect 1610 310 1630 340
rect 980 300 1020 310
rect 980 280 990 300
rect 1010 280 1020 300
rect 980 270 1020 280
rect 1610 300 1650 310
rect 1610 280 1620 300
rect 1640 280 1650 300
rect 1610 270 1650 280
rect 370 240 410 250
rect -40 165 0 175
rect -40 95 -30 165
rect -10 95 0 165
rect -40 85 0 95
rect 110 165 150 175
rect 110 95 120 165
rect 140 95 150 165
rect 110 85 150 95
rect 260 165 300 175
rect 260 95 270 165
rect 290 95 300 165
rect 260 85 300 95
rect -30 -45 -10 85
rect 20 55 60 65
rect 20 35 30 55
rect 50 35 60 55
rect 20 25 60 35
rect -125 -55 -85 -45
rect -125 -125 -115 -55
rect -95 -125 -85 -55
rect -125 -135 -85 -125
rect -40 -55 0 -45
rect -40 -125 -30 -55
rect -10 -125 0 -55
rect -40 -135 0 -125
rect -30 -165 -10 -135
rect 30 -155 50 25
rect 120 -45 140 85
rect 170 55 210 65
rect 170 35 180 55
rect 200 35 210 55
rect 170 25 210 35
rect 270 30 290 85
rect 370 70 380 240
rect 400 70 410 240
rect 370 60 410 70
rect 920 240 960 250
rect 920 70 930 240
rect 950 70 960 240
rect 920 60 960 70
rect 380 30 400 60
rect 110 -55 150 -45
rect 110 -125 120 -55
rect 140 -125 150 -55
rect 110 -135 150 -125
rect 20 -165 60 -155
rect 120 -165 140 -135
rect 180 -155 200 25
rect 270 10 400 30
rect 270 -45 290 10
rect 260 -55 300 -45
rect 260 -125 270 -55
rect 290 -125 300 -55
rect 260 -135 300 -125
rect -30 -185 30 -165
rect 50 -185 140 -165
rect 170 -165 210 -155
rect 170 -185 180 -165
rect 200 -185 210 -165
rect 380 -170 400 10
rect 430 30 470 40
rect 430 10 440 30
rect 460 10 470 30
rect 430 0 470 10
rect 20 -195 60 -185
rect 170 -195 210 -185
rect 370 -180 410 -170
rect 180 -510 200 -195
rect 370 -350 380 -180
rect 400 -350 410 -180
rect 370 -360 410 -350
rect 440 -380 460 0
rect 930 -170 950 60
rect 990 -110 1010 270
rect 1470 240 1510 250
rect 1470 70 1480 240
rect 1500 70 1510 240
rect 1470 60 1510 70
rect 980 -120 1020 -110
rect 980 -140 990 -120
rect 1010 -140 1020 -120
rect 980 -150 1020 -140
rect 1480 -170 1500 60
rect 1535 -20 1575 -10
rect 1535 -90 1545 -20
rect 1565 -90 1575 -20
rect 1535 -100 1575 -90
rect 1620 -110 1640 270
rect 2570 250 2595 340
rect 2020 240 2060 250
rect 2020 70 2030 240
rect 2050 70 2060 240
rect 2020 60 2060 70
rect 2570 240 2610 250
rect 2570 70 2580 240
rect 2600 70 2610 240
rect 2920 140 2940 380
rect 2570 60 2610 70
rect 2760 130 2800 140
rect 2760 60 2770 130
rect 2790 60 2800 130
rect 1610 -120 1650 -110
rect 1610 -140 1620 -120
rect 1640 -140 1650 -120
rect 1610 -150 1650 -140
rect 2030 -170 2050 60
rect 2080 30 2120 40
rect 2080 10 2090 30
rect 2110 10 2120 30
rect 2080 0 2120 10
rect 2580 0 2600 60
rect 2760 50 2800 60
rect 2910 130 2950 140
rect 2910 60 2920 130
rect 2940 60 2950 130
rect 2910 50 2950 60
rect 3060 130 3100 140
rect 3060 60 3070 130
rect 3090 60 3100 130
rect 3060 50 3100 60
rect 2770 0 2790 50
rect 920 -180 960 -170
rect 920 -350 930 -180
rect 950 -350 960 -180
rect 920 -360 960 -350
rect 1470 -180 1510 -170
rect 1470 -350 1480 -180
rect 1500 -350 1510 -180
rect 1470 -360 1510 -350
rect 2020 -180 2060 -170
rect 2020 -350 2030 -180
rect 2050 -350 2060 -180
rect 2020 -360 2060 -350
rect 430 -390 470 -380
rect 430 -410 440 -390
rect 460 -410 470 -390
rect 430 -420 470 -410
rect 930 -395 950 -360
rect 2030 -395 2050 -360
rect 2090 -380 2110 0
rect 2580 -20 2790 0
rect 2820 20 2860 30
rect 2820 0 2830 20
rect 2850 0 2860 20
rect 2820 -10 2860 0
rect 2580 -170 2600 -20
rect 2770 -80 2790 -20
rect 2675 -90 2715 -80
rect 2675 -160 2685 -90
rect 2705 -160 2715 -90
rect 2675 -170 2715 -160
rect 2760 -90 2800 -80
rect 2760 -160 2770 -90
rect 2790 -160 2800 -90
rect 2760 -170 2800 -160
rect 2570 -180 2610 -170
rect 2570 -350 2580 -180
rect 2600 -350 2610 -180
rect 2830 -190 2850 -10
rect 2920 -80 2940 50
rect 2970 20 3010 30
rect 2970 0 2980 20
rect 3000 0 3010 20
rect 2970 -10 3010 0
rect 2910 -90 2950 -80
rect 2910 -160 2920 -90
rect 2940 -160 2950 -90
rect 2910 -170 2950 -160
rect 2570 -360 2610 -350
rect 2820 -200 2860 -190
rect 2820 -220 2830 -200
rect 2850 -220 2860 -200
rect 2920 -200 2940 -170
rect 2980 -190 3000 -10
rect 3070 -80 3090 50
rect 3060 -90 3100 -80
rect 3060 -160 3070 -90
rect 3090 -160 3100 -90
rect 3060 -170 3100 -160
rect 2970 -200 3010 -190
rect 3070 -200 3090 -170
rect 2920 -220 2980 -200
rect 3000 -220 3090 -200
rect 2820 -230 2860 -220
rect 2970 -230 3010 -220
rect 930 -420 2050 -395
rect 2080 -390 2120 -380
rect 2080 -410 2090 -390
rect 2110 -410 2120 -390
rect 2080 -420 2120 -410
rect 440 -460 460 -420
rect 2080 -460 2100 -420
rect 440 -480 2100 -460
rect 2820 -510 2845 -230
rect 180 -530 2845 -510
<< end >>
