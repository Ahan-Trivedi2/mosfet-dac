magic
tech sky130A
timestamp 1762135317
<< nwell >>
rect 4160 6240 4400 7540
rect 7900 6240 8140 7540
rect 4160 4160 8140 6240
rect 4160 2860 4400 4160
rect 7900 2860 8140 4160
<< nmos >>
rect 4460 7520 4560 7620
rect 4630 7520 4730 7620
rect 4800 7520 4900 7620
rect 4970 7520 5070 7620
rect 5140 7520 5240 7620
rect 5310 7520 5410 7620
rect 5480 7520 5580 7620
rect 5650 7520 5750 7620
rect 5820 7520 5920 7620
rect 5990 7520 6090 7620
rect 6210 7520 6310 7620
rect 6380 7520 6480 7620
rect 6550 7520 6650 7620
rect 6720 7520 6820 7620
rect 6890 7520 6990 7620
rect 7060 7520 7160 7620
rect 7230 7520 7330 7620
rect 7400 7520 7500 7620
rect 7570 7520 7670 7620
rect 7740 7520 7840 7620
rect 4460 7380 4560 7480
rect 4630 7380 4730 7480
rect 4800 7380 4900 7480
rect 4970 7380 5070 7480
rect 5140 7380 5240 7480
rect 5310 7380 5410 7480
rect 5480 7380 5580 7480
rect 5650 7380 5750 7480
rect 5820 7380 5920 7480
rect 5990 7380 6090 7480
rect 4460 6340 4560 7340
rect 4630 6340 4730 7340
rect 4800 6340 4900 7340
rect 4970 6340 5070 7340
rect 5140 6340 5240 7340
rect 5310 6340 5410 7340
rect 5480 6340 5580 7340
rect 5650 6340 5750 7340
rect 5820 6340 5920 7340
rect 5990 6340 6090 7340
rect 6210 7380 6310 7480
rect 6380 7380 6480 7480
rect 6550 7380 6650 7480
rect 6720 7380 6820 7480
rect 6890 7380 6990 7480
rect 7060 7380 7160 7480
rect 7230 7380 7330 7480
rect 7400 7380 7500 7480
rect 7570 7380 7670 7480
rect 7740 7380 7840 7480
rect 6210 6340 6310 7340
rect 6380 6340 6480 7340
rect 6550 6340 6650 7340
rect 6720 6340 6820 7340
rect 6890 6340 6990 7340
rect 7060 6340 7160 7340
rect 7230 6340 7330 7340
rect 7400 6340 7500 7340
rect 7570 6340 7670 7340
rect 7740 6340 7840 7340
rect 4460 3060 4560 4060
rect 4630 3060 4730 4060
rect 4800 3060 4900 4060
rect 4970 3060 5070 4060
rect 5140 3060 5240 4060
rect 5310 3060 5410 4060
rect 5480 3060 5580 4060
rect 5650 3060 5750 4060
rect 5820 3060 5920 4060
rect 5990 3060 6090 4060
rect 4460 2920 4560 3020
rect 4630 2920 4730 3020
rect 4800 2920 4900 3020
rect 4970 2920 5070 3020
rect 5140 2920 5240 3020
rect 5310 2920 5410 3020
rect 5480 2920 5580 3020
rect 5650 2920 5750 3020
rect 5820 2920 5920 3020
rect 5990 2920 6090 3020
rect 6210 3060 6310 4060
rect 6380 3060 6480 4060
rect 6550 3060 6650 4060
rect 6720 3060 6820 4060
rect 6890 3060 6990 4060
rect 7060 3060 7160 4060
rect 7230 3060 7330 4060
rect 7400 3060 7500 4060
rect 7570 3060 7670 4060
rect 7740 3060 7840 4060
rect 6210 2920 6310 3020
rect 6380 2920 6480 3020
rect 6550 2920 6650 3020
rect 6720 2920 6820 3020
rect 6890 2920 6990 3020
rect 7060 2920 7160 3020
rect 7230 2920 7330 3020
rect 7400 2920 7500 3020
rect 7570 2920 7670 3020
rect 7740 2920 7840 3020
rect 4460 2780 4560 2880
rect 4630 2780 4730 2880
rect 4800 2780 4900 2880
rect 4970 2780 5070 2880
rect 5140 2780 5240 2880
rect 5310 2780 5410 2880
rect 5480 2780 5580 2880
rect 5650 2780 5750 2880
rect 5820 2780 5920 2880
rect 5990 2780 6090 2880
rect 6210 2780 6310 2880
rect 6380 2780 6480 2880
rect 6550 2780 6650 2880
rect 6720 2780 6820 2880
rect 6890 2780 6990 2880
rect 7060 2780 7160 2880
rect 7230 2780 7330 2880
rect 7400 2780 7500 2880
rect 7570 2780 7670 2880
rect 7740 2780 7840 2880
<< pmos >>
rect 4180 6980 4380 7480
rect 4180 6440 4380 6940
rect 7920 6980 8120 7480
rect 7920 6440 8120 6940
rect 4300 5220 4400 6220
rect 4440 5220 4540 6220
rect 4580 5220 4680 6220
rect 4720 5220 4820 6220
rect 4860 5220 4960 6220
rect 5000 5220 5100 6220
rect 5140 5220 5240 6220
rect 5280 5220 5380 6220
rect 5420 5220 5520 6220
rect 5560 5220 5660 6220
rect 5700 5220 5800 6220
rect 4300 4180 4400 5180
rect 4440 4180 4540 5180
rect 4580 4180 4680 5180
rect 4720 4180 4820 5180
rect 4860 4180 4960 5180
rect 5000 4180 5100 5180
rect 5140 4180 5240 5180
rect 5280 4180 5380 5180
rect 5420 4180 5520 5180
rect 5560 4180 5660 5180
rect 5700 4180 5800 5180
rect 6500 5220 6600 6220
rect 6640 5220 6740 6220
rect 6780 5220 6880 6220
rect 6920 5220 7020 6220
rect 7060 5220 7160 6220
rect 7200 5220 7300 6220
rect 7340 5220 7440 6220
rect 7480 5220 7580 6220
rect 7620 5220 7720 6220
rect 7760 5220 7860 6220
rect 7900 5220 8000 6220
rect 6500 4180 6600 5180
rect 6640 4180 6740 5180
rect 6780 4180 6880 5180
rect 6920 4180 7020 5180
rect 7060 4180 7160 5180
rect 7200 4180 7300 5180
rect 7340 4180 7440 5180
rect 7480 4180 7580 5180
rect 7620 4180 7720 5180
rect 7760 4180 7860 5180
rect 7900 4180 8000 5180
rect 4180 3460 4380 3960
rect 4180 2920 4380 3420
rect 7920 3460 8120 3960
rect 7920 2920 8120 3420
<< ndiff >>
rect 4460 7650 4560 7660
rect 4460 7630 4490 7650
rect 4530 7630 4560 7650
rect 4460 7620 4560 7630
rect 4630 7650 4730 7660
rect 4630 7630 4660 7650
rect 4700 7630 4730 7650
rect 4630 7620 4730 7630
rect 4800 7650 4900 7660
rect 4800 7630 4830 7650
rect 4870 7630 4900 7650
rect 4800 7620 4900 7630
rect 4970 7650 5070 7660
rect 4970 7630 5000 7650
rect 5040 7630 5070 7650
rect 4970 7620 5070 7630
rect 5140 7650 5240 7660
rect 5140 7630 5170 7650
rect 5210 7630 5240 7650
rect 5140 7620 5240 7630
rect 5310 7650 5410 7660
rect 5310 7630 5340 7650
rect 5380 7630 5410 7650
rect 5310 7620 5410 7630
rect 5480 7650 5580 7660
rect 5480 7630 5510 7650
rect 5550 7630 5580 7650
rect 5480 7620 5580 7630
rect 5650 7650 5750 7660
rect 5650 7630 5680 7650
rect 5720 7630 5750 7650
rect 5650 7620 5750 7630
rect 5820 7650 5920 7660
rect 5820 7630 5850 7650
rect 5890 7630 5920 7650
rect 5820 7620 5920 7630
rect 5990 7650 6090 7660
rect 5990 7630 6020 7650
rect 6060 7630 6090 7650
rect 5990 7620 6090 7630
rect 6210 7650 6310 7660
rect 6210 7630 6240 7650
rect 6280 7630 6310 7650
rect 6210 7620 6310 7630
rect 6380 7650 6480 7660
rect 6380 7630 6410 7650
rect 6450 7630 6480 7650
rect 6380 7620 6480 7630
rect 6550 7650 6650 7660
rect 6550 7630 6580 7650
rect 6620 7630 6650 7650
rect 6550 7620 6650 7630
rect 6720 7650 6820 7660
rect 6720 7630 6750 7650
rect 6790 7630 6820 7650
rect 6720 7620 6820 7630
rect 6890 7650 6990 7660
rect 6890 7630 6920 7650
rect 6960 7630 6990 7650
rect 6890 7620 6990 7630
rect 7060 7650 7160 7660
rect 7060 7630 7090 7650
rect 7130 7630 7160 7650
rect 7060 7620 7160 7630
rect 7230 7650 7330 7660
rect 7230 7630 7260 7650
rect 7300 7630 7330 7650
rect 7230 7620 7330 7630
rect 7400 7650 7500 7660
rect 7400 7630 7430 7650
rect 7470 7630 7500 7650
rect 7400 7620 7500 7630
rect 7570 7650 7670 7660
rect 7570 7630 7600 7650
rect 7640 7630 7670 7650
rect 7570 7620 7670 7630
rect 7740 7650 7840 7660
rect 7740 7630 7770 7650
rect 7810 7630 7840 7650
rect 7740 7620 7840 7630
rect 4460 7510 4560 7520
rect 4630 7510 4730 7520
rect 4800 7510 4900 7520
rect 4970 7510 5070 7520
rect 5140 7510 5240 7520
rect 5310 7510 5410 7520
rect 5480 7510 5580 7520
rect 5650 7510 5750 7520
rect 5820 7510 5920 7520
rect 5990 7510 6090 7520
rect 6210 7510 6310 7520
rect 6380 7510 6480 7520
rect 6550 7510 6650 7520
rect 6720 7510 6820 7520
rect 6890 7510 6990 7520
rect 7060 7510 7160 7520
rect 7230 7510 7330 7520
rect 7400 7510 7500 7520
rect 7570 7510 7670 7520
rect 7740 7510 7840 7520
rect 4460 7490 4490 7510
rect 4530 7490 4660 7510
rect 4700 7490 4830 7510
rect 4870 7490 5000 7510
rect 5040 7490 5170 7510
rect 5210 7490 5340 7510
rect 5380 7490 5510 7510
rect 5550 7490 5680 7510
rect 5720 7490 5850 7510
rect 5890 7490 6020 7510
rect 6060 7490 6240 7510
rect 6280 7490 6410 7510
rect 6450 7490 6580 7510
rect 6620 7490 6750 7510
rect 6790 7490 6920 7510
rect 6960 7490 7090 7510
rect 7130 7490 7260 7510
rect 7300 7490 7430 7510
rect 7470 7490 7600 7510
rect 7640 7490 7770 7510
rect 7810 7490 7840 7510
rect 4460 7480 4560 7490
rect 4630 7480 4730 7490
rect 4800 7480 4900 7490
rect 4970 7480 5070 7490
rect 5140 7480 5240 7490
rect 5310 7480 5410 7490
rect 5480 7480 5580 7490
rect 5650 7480 5750 7490
rect 5820 7480 5920 7490
rect 5990 7480 6090 7490
rect 6210 7480 6310 7490
rect 6380 7480 6480 7490
rect 6550 7480 6650 7490
rect 6720 7480 6820 7490
rect 6890 7480 6990 7490
rect 7060 7480 7160 7490
rect 7230 7480 7330 7490
rect 7400 7480 7500 7490
rect 7570 7480 7670 7490
rect 7740 7480 7840 7490
rect 4460 7370 4560 7380
rect 4460 7350 4490 7370
rect 4530 7350 4560 7370
rect 4460 7340 4560 7350
rect 4630 7370 4730 7380
rect 4630 7350 4660 7370
rect 4700 7350 4730 7370
rect 4630 7340 4730 7350
rect 4800 7370 4900 7380
rect 4800 7350 4830 7370
rect 4870 7350 4900 7370
rect 4800 7340 4900 7350
rect 4970 7370 5070 7380
rect 4970 7350 5000 7370
rect 5040 7350 5070 7370
rect 4970 7340 5070 7350
rect 5140 7370 5240 7380
rect 5140 7350 5170 7370
rect 5210 7350 5240 7370
rect 5140 7340 5240 7350
rect 5310 7370 5410 7380
rect 5310 7350 5340 7370
rect 5380 7350 5410 7370
rect 5310 7340 5410 7350
rect 5480 7370 5580 7380
rect 5480 7350 5510 7370
rect 5550 7350 5580 7370
rect 5480 7340 5580 7350
rect 5650 7370 5750 7380
rect 5650 7350 5680 7370
rect 5720 7350 5750 7370
rect 5650 7340 5750 7350
rect 5820 7370 5920 7380
rect 5820 7350 5850 7370
rect 5890 7350 5920 7370
rect 5820 7340 5920 7350
rect 5990 7370 6090 7380
rect 5990 7350 6020 7370
rect 6060 7350 6090 7370
rect 5990 7340 6090 7350
rect 6210 7370 6310 7380
rect 6210 7350 6240 7370
rect 6280 7350 6310 7370
rect 6210 7340 6310 7350
rect 6380 7370 6480 7380
rect 6380 7350 6410 7370
rect 6450 7350 6480 7370
rect 6380 7340 6480 7350
rect 6550 7370 6650 7380
rect 6550 7350 6580 7370
rect 6620 7350 6650 7370
rect 6550 7340 6650 7350
rect 6720 7370 6820 7380
rect 6720 7350 6750 7370
rect 6790 7350 6820 7370
rect 6720 7340 6820 7350
rect 6890 7370 6990 7380
rect 6890 7350 6920 7370
rect 6960 7350 6990 7370
rect 6890 7340 6990 7350
rect 7060 7370 7160 7380
rect 7060 7350 7090 7370
rect 7130 7350 7160 7370
rect 7060 7340 7160 7350
rect 7230 7370 7330 7380
rect 7230 7350 7260 7370
rect 7300 7350 7330 7370
rect 7230 7340 7330 7350
rect 7400 7370 7500 7380
rect 7400 7350 7430 7370
rect 7470 7350 7500 7370
rect 7400 7340 7500 7350
rect 7570 7370 7670 7380
rect 7570 7350 7600 7370
rect 7640 7350 7670 7370
rect 7570 7340 7670 7350
rect 7740 7370 7840 7380
rect 7740 7350 7770 7370
rect 7810 7350 7840 7370
rect 7740 7340 7840 7350
rect 4460 6330 4560 6340
rect 4460 6310 4490 6330
rect 4530 6310 4560 6330
rect 4460 6300 4560 6310
rect 4630 6330 4730 6340
rect 4630 6310 4660 6330
rect 4700 6310 4730 6330
rect 4630 6300 4730 6310
rect 4800 6330 4900 6340
rect 4800 6310 4830 6330
rect 4870 6310 4900 6330
rect 4800 6300 4900 6310
rect 4970 6330 5070 6340
rect 4970 6310 5000 6330
rect 5040 6310 5070 6330
rect 4970 6300 5070 6310
rect 5140 6330 5240 6340
rect 5140 6310 5170 6330
rect 5210 6310 5240 6330
rect 5140 6300 5240 6310
rect 5310 6330 5410 6340
rect 5310 6310 5340 6330
rect 5380 6310 5410 6330
rect 5310 6300 5410 6310
rect 5480 6330 5580 6340
rect 5480 6310 5510 6330
rect 5550 6310 5580 6330
rect 5480 6300 5580 6310
rect 5650 6330 5750 6340
rect 5650 6310 5680 6330
rect 5720 6310 5750 6330
rect 5650 6300 5750 6310
rect 5820 6330 5920 6340
rect 5820 6310 5850 6330
rect 5890 6310 5920 6330
rect 5820 6300 5920 6310
rect 5990 6330 6090 6340
rect 5990 6310 6020 6330
rect 6060 6310 6090 6330
rect 5990 6300 6090 6310
rect 6210 6330 6310 6340
rect 6210 6310 6240 6330
rect 6280 6310 6310 6330
rect 6210 6300 6310 6310
rect 6380 6330 6480 6340
rect 6380 6310 6410 6330
rect 6450 6310 6480 6330
rect 6380 6300 6480 6310
rect 6550 6330 6650 6340
rect 6550 6310 6580 6330
rect 6620 6310 6650 6330
rect 6550 6300 6650 6310
rect 6720 6330 6820 6340
rect 6720 6310 6750 6330
rect 6790 6310 6820 6330
rect 6720 6300 6820 6310
rect 6890 6330 6990 6340
rect 6890 6310 6920 6330
rect 6960 6310 6990 6330
rect 6890 6300 6990 6310
rect 7060 6330 7160 6340
rect 7060 6310 7090 6330
rect 7130 6310 7160 6330
rect 7060 6300 7160 6310
rect 7230 6330 7330 6340
rect 7230 6310 7260 6330
rect 7300 6310 7330 6330
rect 7230 6300 7330 6310
rect 7400 6330 7500 6340
rect 7400 6310 7430 6330
rect 7470 6310 7500 6330
rect 7400 6300 7500 6310
rect 7570 6330 7670 6340
rect 7570 6310 7600 6330
rect 7640 6310 7670 6330
rect 7570 6300 7670 6310
rect 7740 6330 7840 6340
rect 7740 6310 7770 6330
rect 7810 6310 7840 6330
rect 7740 6300 7840 6310
rect 4460 4090 4560 4100
rect 4460 4070 4490 4090
rect 4530 4070 4560 4090
rect 4460 4060 4560 4070
rect 4630 4090 4730 4100
rect 4630 4070 4660 4090
rect 4700 4070 4730 4090
rect 4630 4060 4730 4070
rect 4800 4090 4900 4100
rect 4800 4070 4830 4090
rect 4870 4070 4900 4090
rect 4800 4060 4900 4070
rect 4970 4090 5070 4100
rect 4970 4070 5000 4090
rect 5040 4070 5070 4090
rect 4970 4060 5070 4070
rect 5140 4090 5240 4100
rect 5140 4070 5170 4090
rect 5210 4070 5240 4090
rect 5140 4060 5240 4070
rect 5310 4090 5410 4100
rect 5310 4070 5340 4090
rect 5380 4070 5410 4090
rect 5310 4060 5410 4070
rect 5480 4090 5580 4100
rect 5480 4070 5510 4090
rect 5550 4070 5580 4090
rect 5480 4060 5580 4070
rect 5650 4090 5750 4100
rect 5650 4070 5680 4090
rect 5720 4070 5750 4090
rect 5650 4060 5750 4070
rect 5820 4090 5920 4100
rect 5820 4070 5850 4090
rect 5890 4070 5920 4090
rect 5820 4060 5920 4070
rect 5990 4090 6090 4100
rect 5990 4070 6020 4090
rect 6060 4070 6090 4090
rect 5990 4060 6090 4070
rect 6210 4090 6310 4100
rect 6210 4070 6240 4090
rect 6280 4070 6310 4090
rect 6210 4060 6310 4070
rect 6380 4090 6480 4100
rect 6380 4070 6410 4090
rect 6450 4070 6480 4090
rect 6380 4060 6480 4070
rect 6550 4090 6650 4100
rect 6550 4070 6580 4090
rect 6620 4070 6650 4090
rect 6550 4060 6650 4070
rect 6720 4090 6820 4100
rect 6720 4070 6750 4090
rect 6790 4070 6820 4090
rect 6720 4060 6820 4070
rect 6890 4090 6990 4100
rect 6890 4070 6920 4090
rect 6960 4070 6990 4090
rect 6890 4060 6990 4070
rect 7060 4090 7160 4100
rect 7060 4070 7090 4090
rect 7130 4070 7160 4090
rect 7060 4060 7160 4070
rect 7230 4090 7330 4100
rect 7230 4070 7260 4090
rect 7300 4070 7330 4090
rect 7230 4060 7330 4070
rect 7400 4090 7500 4100
rect 7400 4070 7430 4090
rect 7470 4070 7500 4090
rect 7400 4060 7500 4070
rect 7570 4090 7670 4100
rect 7570 4070 7600 4090
rect 7640 4070 7670 4090
rect 7570 4060 7670 4070
rect 7740 4090 7840 4100
rect 7740 4070 7770 4090
rect 7810 4070 7840 4090
rect 7740 4060 7840 4070
rect 4460 3050 4560 3060
rect 4460 3030 4490 3050
rect 4530 3030 4560 3050
rect 4460 3020 4560 3030
rect 4630 3050 4730 3060
rect 4630 3030 4660 3050
rect 4700 3030 4730 3050
rect 4630 3020 4730 3030
rect 4800 3050 4900 3060
rect 4800 3030 4830 3050
rect 4870 3030 4900 3050
rect 4800 3020 4900 3030
rect 4970 3050 5070 3060
rect 4970 3030 5000 3050
rect 5040 3030 5070 3050
rect 4970 3020 5070 3030
rect 5140 3050 5240 3060
rect 5140 3030 5170 3050
rect 5210 3030 5240 3050
rect 5140 3020 5240 3030
rect 5310 3050 5410 3060
rect 5310 3030 5340 3050
rect 5380 3030 5410 3050
rect 5310 3020 5410 3030
rect 5480 3050 5580 3060
rect 5480 3030 5510 3050
rect 5550 3030 5580 3050
rect 5480 3020 5580 3030
rect 5650 3050 5750 3060
rect 5650 3030 5680 3050
rect 5720 3030 5750 3050
rect 5650 3020 5750 3030
rect 5820 3050 5920 3060
rect 5820 3030 5850 3050
rect 5890 3030 5920 3050
rect 5820 3020 5920 3030
rect 5990 3050 6090 3060
rect 5990 3030 6020 3050
rect 6060 3030 6090 3050
rect 5990 3020 6090 3030
rect 6210 3050 6310 3060
rect 6210 3030 6240 3050
rect 6280 3030 6310 3050
rect 6210 3020 6310 3030
rect 6380 3050 6480 3060
rect 6380 3030 6410 3050
rect 6450 3030 6480 3050
rect 6380 3020 6480 3030
rect 6550 3050 6650 3060
rect 6550 3030 6580 3050
rect 6620 3030 6650 3050
rect 6550 3020 6650 3030
rect 6720 3050 6820 3060
rect 6720 3030 6750 3050
rect 6790 3030 6820 3050
rect 6720 3020 6820 3030
rect 6890 3050 6990 3060
rect 6890 3030 6920 3050
rect 6960 3030 6990 3050
rect 6890 3020 6990 3030
rect 7060 3050 7160 3060
rect 7060 3030 7090 3050
rect 7130 3030 7160 3050
rect 7060 3020 7160 3030
rect 7230 3050 7330 3060
rect 7230 3030 7260 3050
rect 7300 3030 7330 3050
rect 7230 3020 7330 3030
rect 7400 3050 7500 3060
rect 7400 3030 7430 3050
rect 7470 3030 7500 3050
rect 7400 3020 7500 3030
rect 7570 3050 7670 3060
rect 7570 3030 7600 3050
rect 7640 3030 7670 3050
rect 7570 3020 7670 3030
rect 7740 3050 7840 3060
rect 7740 3030 7770 3050
rect 7810 3030 7840 3050
rect 7740 3020 7840 3030
rect 4460 2910 4560 2920
rect 4630 2910 4730 2920
rect 4800 2910 4900 2920
rect 4970 2910 5070 2920
rect 5140 2910 5240 2920
rect 5310 2910 5410 2920
rect 5480 2910 5580 2920
rect 5650 2910 5750 2920
rect 5820 2910 5920 2920
rect 5990 2910 6090 2920
rect 6210 2910 6310 2920
rect 6380 2910 6480 2920
rect 6550 2910 6650 2920
rect 6720 2910 6820 2920
rect 6890 2910 6990 2920
rect 7060 2910 7160 2920
rect 7230 2910 7330 2920
rect 7400 2910 7500 2920
rect 7570 2910 7670 2920
rect 7740 2910 7840 2920
rect 4460 2890 4490 2910
rect 4530 2890 4660 2910
rect 4700 2890 4830 2910
rect 4870 2890 5000 2910
rect 5040 2890 5170 2910
rect 5210 2890 5340 2910
rect 5380 2890 5510 2910
rect 5550 2890 5680 2910
rect 5720 2890 5850 2910
rect 5890 2890 6020 2910
rect 6060 2890 6240 2910
rect 6280 2890 6410 2910
rect 6450 2890 6580 2910
rect 6620 2890 6750 2910
rect 6790 2890 6920 2910
rect 6960 2890 7090 2910
rect 7130 2890 7260 2910
rect 7300 2890 7430 2910
rect 7470 2890 7600 2910
rect 7640 2890 7770 2910
rect 7810 2890 7840 2910
rect 4460 2880 4560 2890
rect 4630 2880 4730 2890
rect 4800 2880 4900 2890
rect 4970 2880 5070 2890
rect 5140 2880 5240 2890
rect 5310 2880 5410 2890
rect 5480 2880 5580 2890
rect 5650 2880 5750 2890
rect 5820 2880 5920 2890
rect 5990 2880 6090 2890
rect 6210 2880 6310 2890
rect 6380 2880 6480 2890
rect 6550 2880 6650 2890
rect 6720 2880 6820 2890
rect 6890 2880 6990 2890
rect 7060 2880 7160 2890
rect 7230 2880 7330 2890
rect 7400 2880 7500 2890
rect 7570 2880 7670 2890
rect 7740 2880 7840 2890
rect 4460 2770 4560 2780
rect 4460 2750 4490 2770
rect 4530 2750 4560 2770
rect 4460 2740 4560 2750
rect 4630 2770 4730 2780
rect 4630 2750 4660 2770
rect 4700 2750 4730 2770
rect 4630 2740 4730 2750
rect 4800 2770 4900 2780
rect 4800 2750 4830 2770
rect 4870 2750 4900 2770
rect 4800 2740 4900 2750
rect 4970 2770 5070 2780
rect 4970 2750 5000 2770
rect 5040 2750 5070 2770
rect 4970 2740 5070 2750
rect 5140 2770 5240 2780
rect 5140 2750 5170 2770
rect 5210 2750 5240 2770
rect 5140 2740 5240 2750
rect 5310 2770 5410 2780
rect 5310 2750 5340 2770
rect 5380 2750 5410 2770
rect 5310 2740 5410 2750
rect 5480 2770 5580 2780
rect 5480 2750 5510 2770
rect 5550 2750 5580 2770
rect 5480 2740 5580 2750
rect 5650 2770 5750 2780
rect 5650 2750 5680 2770
rect 5720 2750 5750 2770
rect 5650 2740 5750 2750
rect 5820 2770 5920 2780
rect 5820 2750 5850 2770
rect 5890 2750 5920 2770
rect 5820 2740 5920 2750
rect 5990 2770 6090 2780
rect 5990 2750 6020 2770
rect 6060 2750 6090 2770
rect 5990 2740 6090 2750
rect 6210 2770 6310 2780
rect 6210 2750 6240 2770
rect 6280 2750 6310 2770
rect 6210 2740 6310 2750
rect 6380 2770 6480 2780
rect 6380 2750 6410 2770
rect 6450 2750 6480 2770
rect 6380 2740 6480 2750
rect 6550 2770 6650 2780
rect 6550 2750 6580 2770
rect 6620 2750 6650 2770
rect 6550 2740 6650 2750
rect 6720 2770 6820 2780
rect 6720 2750 6750 2770
rect 6790 2750 6820 2770
rect 6720 2740 6820 2750
rect 6890 2770 6990 2780
rect 6890 2750 6920 2770
rect 6960 2750 6990 2770
rect 6890 2740 6990 2750
rect 7060 2770 7160 2780
rect 7060 2750 7090 2770
rect 7130 2750 7160 2770
rect 7060 2740 7160 2750
rect 7230 2770 7330 2780
rect 7230 2750 7260 2770
rect 7300 2750 7330 2770
rect 7230 2740 7330 2750
rect 7400 2770 7500 2780
rect 7400 2750 7430 2770
rect 7470 2750 7500 2770
rect 7400 2740 7500 2750
rect 7570 2770 7670 2780
rect 7570 2750 7600 2770
rect 7640 2750 7670 2770
rect 7570 2740 7670 2750
rect 7740 2770 7840 2780
rect 7740 2750 7770 2770
rect 7810 2750 7840 2770
rect 7740 2740 7840 2750
<< pdiff >>
rect 4180 7510 4380 7520
rect 4180 7490 4260 7510
rect 4300 7490 4380 7510
rect 4180 7480 4380 7490
rect 7920 7510 8120 7520
rect 7920 7490 8000 7510
rect 8040 7490 8120 7510
rect 7920 7480 8120 7490
rect 4180 6970 4380 6980
rect 4180 6950 4260 6970
rect 4300 6950 4380 6970
rect 4180 6940 4380 6950
rect 4180 6430 4380 6440
rect 4180 6410 4240 6430
rect 4280 6410 4380 6430
rect 4180 6400 4380 6410
rect 7920 6970 8120 6980
rect 7920 6950 8000 6970
rect 8040 6950 8120 6970
rect 7920 6940 8120 6950
rect 7920 6430 8120 6440
rect 7920 6410 8020 6430
rect 8060 6410 8120 6430
rect 7920 6400 8120 6410
rect 4220 6200 4300 6220
rect 4260 6140 4300 6200
rect 4220 5740 4300 6140
rect 4220 5700 4270 5740
rect 4290 5700 4300 5740
rect 4220 5220 4300 5700
rect 4400 5740 4440 6220
rect 4400 5700 4410 5740
rect 4430 5700 4440 5740
rect 4400 5220 4440 5700
rect 4540 5740 4580 6220
rect 4540 5700 4550 5740
rect 4570 5700 4580 5740
rect 4540 5220 4580 5700
rect 4680 5740 4720 6220
rect 4680 5700 4690 5740
rect 4710 5700 4720 5740
rect 4680 5220 4720 5700
rect 4820 5740 4860 6220
rect 4820 5700 4830 5740
rect 4850 5700 4860 5740
rect 4820 5220 4860 5700
rect 4960 5740 5000 6220
rect 4960 5700 4970 5740
rect 4990 5700 5000 5740
rect 4960 5220 5000 5700
rect 5100 5740 5140 6220
rect 5100 5700 5110 5740
rect 5130 5700 5140 5740
rect 5100 5220 5140 5700
rect 5240 5740 5280 6220
rect 5240 5700 5250 5740
rect 5270 5700 5280 5740
rect 5240 5220 5280 5700
rect 5380 5740 5420 6220
rect 5380 5700 5390 5740
rect 5410 5700 5420 5740
rect 5380 5220 5420 5700
rect 5520 5740 5560 6220
rect 5520 5700 5530 5740
rect 5550 5700 5560 5740
rect 5520 5220 5560 5700
rect 5660 5740 5700 6220
rect 5660 5700 5670 5740
rect 5690 5700 5700 5740
rect 5660 5220 5700 5700
rect 5800 5740 5840 6220
rect 6010 6210 6290 6220
rect 6010 6190 6020 6210
rect 6040 6190 6260 6210
rect 6280 6190 6290 6210
rect 6010 6180 6290 6190
rect 6460 5740 6500 6220
rect 5800 5700 5810 5740
rect 5830 5700 5840 5740
rect 6010 5730 6290 5740
rect 6010 5710 6020 5730
rect 6040 5710 6260 5730
rect 6280 5710 6290 5730
rect 6010 5700 6290 5710
rect 6460 5700 6470 5740
rect 6490 5700 6500 5740
rect 5800 5220 5840 5700
rect 4220 5180 4290 5220
rect 4410 5180 4430 5220
rect 4550 5180 4570 5220
rect 4690 5180 4710 5220
rect 4830 5180 4850 5220
rect 4970 5180 4990 5220
rect 5110 5180 5130 5220
rect 5250 5180 5270 5220
rect 5390 5180 5410 5220
rect 5530 5180 5550 5220
rect 5670 5180 5690 5220
rect 5810 5180 5830 5220
rect 4220 4700 4300 5180
rect 4220 4660 4270 4700
rect 4290 4660 4300 4700
rect 4220 4260 4300 4660
rect 4260 4200 4300 4260
rect 4220 4180 4300 4200
rect 4400 4700 4440 5180
rect 4400 4660 4410 4700
rect 4430 4660 4440 4700
rect 4400 4180 4440 4660
rect 4540 4700 4580 5180
rect 4540 4660 4550 4700
rect 4570 4660 4580 4700
rect 4540 4180 4580 4660
rect 4680 4700 4720 5180
rect 4680 4660 4690 4700
rect 4710 4660 4720 4700
rect 4680 4180 4720 4660
rect 4820 4700 4860 5180
rect 4820 4660 4830 4700
rect 4850 4660 4860 4700
rect 4820 4180 4860 4660
rect 4960 4700 5000 5180
rect 4960 4660 4970 4700
rect 4990 4660 5000 4700
rect 4960 4180 5000 4660
rect 5100 4700 5140 5180
rect 5100 4660 5110 4700
rect 5130 4660 5140 4700
rect 5100 4180 5140 4660
rect 5240 4700 5280 5180
rect 5240 4660 5250 4700
rect 5270 4660 5280 4700
rect 5240 4180 5280 4660
rect 5380 4700 5420 5180
rect 5380 4660 5390 4700
rect 5410 4660 5420 4700
rect 5380 4180 5420 4660
rect 5520 4700 5560 5180
rect 5520 4660 5530 4700
rect 5550 4660 5560 4700
rect 5520 4180 5560 4660
rect 5660 4700 5700 5180
rect 5660 4660 5670 4700
rect 5690 4660 5700 4700
rect 5660 4180 5700 4660
rect 5800 4700 5840 5180
rect 6010 5210 6290 5220
rect 6010 5190 6020 5210
rect 6040 5190 6260 5210
rect 6280 5190 6290 5210
rect 6010 5180 6290 5190
rect 6460 5220 6500 5700
rect 6600 5740 6640 6220
rect 6600 5700 6610 5740
rect 6630 5700 6640 5740
rect 6600 5220 6640 5700
rect 6740 5740 6780 6220
rect 6740 5700 6750 5740
rect 6770 5700 6780 5740
rect 6740 5220 6780 5700
rect 6880 5740 6920 6220
rect 6880 5700 6890 5740
rect 6910 5700 6920 5740
rect 6880 5220 6920 5700
rect 7020 5740 7060 6220
rect 7020 5700 7030 5740
rect 7050 5700 7060 5740
rect 7020 5220 7060 5700
rect 7160 5740 7200 6220
rect 7160 5700 7170 5740
rect 7190 5700 7200 5740
rect 7160 5220 7200 5700
rect 7300 5740 7340 6220
rect 7300 5700 7310 5740
rect 7330 5700 7340 5740
rect 7300 5220 7340 5700
rect 7440 5740 7480 6220
rect 7440 5700 7450 5740
rect 7470 5700 7480 5740
rect 7440 5220 7480 5700
rect 7580 5740 7620 6220
rect 7580 5700 7590 5740
rect 7610 5700 7620 5740
rect 7580 5220 7620 5700
rect 7720 5740 7760 6220
rect 7720 5700 7730 5740
rect 7750 5700 7760 5740
rect 7720 5220 7760 5700
rect 7860 5740 7900 6220
rect 7860 5700 7870 5740
rect 7890 5700 7900 5740
rect 7860 5220 7900 5700
rect 8000 6200 8080 6220
rect 8000 6140 8040 6200
rect 8000 5740 8080 6140
rect 8000 5700 8010 5740
rect 8030 5700 8080 5740
rect 8000 5220 8080 5700
rect 6470 5180 6490 5220
rect 6610 5180 6630 5220
rect 6750 5180 6770 5220
rect 6890 5180 6910 5220
rect 7030 5180 7050 5220
rect 7170 5180 7190 5220
rect 7310 5180 7330 5220
rect 7450 5180 7470 5220
rect 7590 5180 7610 5220
rect 7730 5180 7750 5220
rect 7870 5180 7890 5220
rect 8010 5180 8080 5220
rect 6460 4700 6500 5180
rect 5800 4660 5810 4700
rect 5830 4660 5840 4700
rect 6010 4690 6290 4700
rect 6010 4670 6020 4690
rect 6040 4670 6260 4690
rect 6280 4670 6290 4690
rect 6010 4660 6290 4670
rect 6460 4660 6470 4700
rect 6490 4660 6500 4700
rect 5800 4180 5840 4660
rect 6010 4210 6290 4220
rect 6010 4190 6020 4210
rect 6040 4190 6260 4210
rect 6280 4190 6290 4210
rect 6010 4180 6290 4190
rect 6460 4180 6500 4660
rect 6600 4700 6640 5180
rect 6600 4660 6610 4700
rect 6630 4660 6640 4700
rect 6600 4180 6640 4660
rect 6740 4700 6780 5180
rect 6740 4660 6750 4700
rect 6770 4660 6780 4700
rect 6740 4180 6780 4660
rect 6880 4700 6920 5180
rect 6880 4660 6890 4700
rect 6910 4660 6920 4700
rect 6880 4180 6920 4660
rect 7020 4700 7060 5180
rect 7020 4660 7030 4700
rect 7050 4660 7060 4700
rect 7020 4180 7060 4660
rect 7160 4700 7200 5180
rect 7160 4660 7170 4700
rect 7190 4660 7200 4700
rect 7160 4180 7200 4660
rect 7300 4700 7340 5180
rect 7300 4660 7310 4700
rect 7330 4660 7340 4700
rect 7300 4180 7340 4660
rect 7440 4700 7480 5180
rect 7440 4660 7450 4700
rect 7470 4660 7480 4700
rect 7440 4180 7480 4660
rect 7580 4700 7620 5180
rect 7580 4660 7590 4700
rect 7610 4660 7620 4700
rect 7580 4180 7620 4660
rect 7720 4700 7760 5180
rect 7720 4660 7730 4700
rect 7750 4660 7760 4700
rect 7720 4180 7760 4660
rect 7860 4700 7900 5180
rect 7860 4660 7870 4700
rect 7890 4660 7900 4700
rect 7860 4180 7900 4660
rect 8000 4700 8080 5180
rect 8000 4660 8010 4700
rect 8030 4660 8080 4700
rect 8000 4260 8080 4660
rect 8000 4200 8040 4260
rect 8000 4180 8080 4200
rect 4180 3990 4380 4000
rect 4180 3970 4240 3990
rect 4280 3970 4380 3990
rect 4180 3960 4380 3970
rect 4180 3450 4380 3460
rect 4180 3430 4260 3450
rect 4300 3430 4380 3450
rect 4180 3420 4380 3430
rect 7920 3990 8120 4000
rect 7920 3970 8020 3990
rect 8060 3970 8120 3990
rect 7920 3960 8120 3970
rect 7920 3450 8120 3460
rect 7920 3430 8000 3450
rect 8040 3430 8120 3450
rect 7920 3420 8120 3430
rect 4180 2910 4380 2920
rect 4180 2890 4260 2910
rect 4300 2890 4380 2910
rect 4180 2880 4380 2890
rect 7920 2910 8120 2920
rect 7920 2890 8000 2910
rect 8040 2890 8120 2910
rect 7920 2880 8120 2890
<< ndiffc >>
rect 4490 7630 4530 7650
rect 4660 7630 4700 7650
rect 4830 7630 4870 7650
rect 5000 7630 5040 7650
rect 5170 7630 5210 7650
rect 5340 7630 5380 7650
rect 5510 7630 5550 7650
rect 5680 7630 5720 7650
rect 5850 7630 5890 7650
rect 6020 7630 6060 7650
rect 6240 7630 6280 7650
rect 6410 7630 6450 7650
rect 6580 7630 6620 7650
rect 6750 7630 6790 7650
rect 6920 7630 6960 7650
rect 7090 7630 7130 7650
rect 7260 7630 7300 7650
rect 7430 7630 7470 7650
rect 7600 7630 7640 7650
rect 7770 7630 7810 7650
rect 4490 7490 4530 7510
rect 4660 7490 4700 7510
rect 4830 7490 4870 7510
rect 5000 7490 5040 7510
rect 5170 7490 5210 7510
rect 5340 7490 5380 7510
rect 5510 7490 5550 7510
rect 5680 7490 5720 7510
rect 5850 7490 5890 7510
rect 6020 7490 6060 7510
rect 6240 7490 6280 7510
rect 6410 7490 6450 7510
rect 6580 7490 6620 7510
rect 6750 7490 6790 7510
rect 6920 7490 6960 7510
rect 7090 7490 7130 7510
rect 7260 7490 7300 7510
rect 7430 7490 7470 7510
rect 7600 7490 7640 7510
rect 7770 7490 7810 7510
rect 4490 7350 4530 7370
rect 4660 7350 4700 7370
rect 4830 7350 4870 7370
rect 5000 7350 5040 7370
rect 5170 7350 5210 7370
rect 5340 7350 5380 7370
rect 5510 7350 5550 7370
rect 5680 7350 5720 7370
rect 5850 7350 5890 7370
rect 6020 7350 6060 7370
rect 6240 7350 6280 7370
rect 6410 7350 6450 7370
rect 6580 7350 6620 7370
rect 6750 7350 6790 7370
rect 6920 7350 6960 7370
rect 7090 7350 7130 7370
rect 7260 7350 7300 7370
rect 7430 7350 7470 7370
rect 7600 7350 7640 7370
rect 7770 7350 7810 7370
rect 4490 6310 4530 6330
rect 4660 6310 4700 6330
rect 4830 6310 4870 6330
rect 5000 6310 5040 6330
rect 5170 6310 5210 6330
rect 5340 6310 5380 6330
rect 5510 6310 5550 6330
rect 5680 6310 5720 6330
rect 5850 6310 5890 6330
rect 6020 6310 6060 6330
rect 6240 6310 6280 6330
rect 6410 6310 6450 6330
rect 6580 6310 6620 6330
rect 6750 6310 6790 6330
rect 6920 6310 6960 6330
rect 7090 6310 7130 6330
rect 7260 6310 7300 6330
rect 7430 6310 7470 6330
rect 7600 6310 7640 6330
rect 7770 6310 7810 6330
rect 4490 4070 4530 4090
rect 4660 4070 4700 4090
rect 4830 4070 4870 4090
rect 5000 4070 5040 4090
rect 5170 4070 5210 4090
rect 5340 4070 5380 4090
rect 5510 4070 5550 4090
rect 5680 4070 5720 4090
rect 5850 4070 5890 4090
rect 6020 4070 6060 4090
rect 6240 4070 6280 4090
rect 6410 4070 6450 4090
rect 6580 4070 6620 4090
rect 6750 4070 6790 4090
rect 6920 4070 6960 4090
rect 7090 4070 7130 4090
rect 7260 4070 7300 4090
rect 7430 4070 7470 4090
rect 7600 4070 7640 4090
rect 7770 4070 7810 4090
rect 4490 3030 4530 3050
rect 4660 3030 4700 3050
rect 4830 3030 4870 3050
rect 5000 3030 5040 3050
rect 5170 3030 5210 3050
rect 5340 3030 5380 3050
rect 5510 3030 5550 3050
rect 5680 3030 5720 3050
rect 5850 3030 5890 3050
rect 6020 3030 6060 3050
rect 6240 3030 6280 3050
rect 6410 3030 6450 3050
rect 6580 3030 6620 3050
rect 6750 3030 6790 3050
rect 6920 3030 6960 3050
rect 7090 3030 7130 3050
rect 7260 3030 7300 3050
rect 7430 3030 7470 3050
rect 7600 3030 7640 3050
rect 7770 3030 7810 3050
rect 4490 2890 4530 2910
rect 4660 2890 4700 2910
rect 4830 2890 4870 2910
rect 5000 2890 5040 2910
rect 5170 2890 5210 2910
rect 5340 2890 5380 2910
rect 5510 2890 5550 2910
rect 5680 2890 5720 2910
rect 5850 2890 5890 2910
rect 6020 2890 6060 2910
rect 6240 2890 6280 2910
rect 6410 2890 6450 2910
rect 6580 2890 6620 2910
rect 6750 2890 6790 2910
rect 6920 2890 6960 2910
rect 7090 2890 7130 2910
rect 7260 2890 7300 2910
rect 7430 2890 7470 2910
rect 7600 2890 7640 2910
rect 7770 2890 7810 2910
rect 4490 2750 4530 2770
rect 4660 2750 4700 2770
rect 4830 2750 4870 2770
rect 5000 2750 5040 2770
rect 5170 2750 5210 2770
rect 5340 2750 5380 2770
rect 5510 2750 5550 2770
rect 5680 2750 5720 2770
rect 5850 2750 5890 2770
rect 6020 2750 6060 2770
rect 6240 2750 6280 2770
rect 6410 2750 6450 2770
rect 6580 2750 6620 2770
rect 6750 2750 6790 2770
rect 6920 2750 6960 2770
rect 7090 2750 7130 2770
rect 7260 2750 7300 2770
rect 7430 2750 7470 2770
rect 7600 2750 7640 2770
rect 7770 2750 7810 2770
<< pdiffc >>
rect 4260 7490 4300 7510
rect 8000 7490 8040 7510
rect 4260 6950 4300 6970
rect 4240 6410 4280 6430
rect 8000 6950 8040 6970
rect 8020 6410 8060 6430
rect 4270 5700 4290 5740
rect 4410 5700 4430 5740
rect 4550 5700 4570 5740
rect 4690 5700 4710 5740
rect 4830 5700 4850 5740
rect 4970 5700 4990 5740
rect 5110 5700 5130 5740
rect 5250 5700 5270 5740
rect 5390 5700 5410 5740
rect 5530 5700 5550 5740
rect 5670 5700 5690 5740
rect 6020 6190 6040 6210
rect 6260 6190 6280 6210
rect 5810 5700 5830 5740
rect 6020 5710 6040 5730
rect 6260 5710 6280 5730
rect 6470 5700 6490 5740
rect 4270 4660 4290 4700
rect 4410 4660 4430 4700
rect 4550 4660 4570 4700
rect 4690 4660 4710 4700
rect 4830 4660 4850 4700
rect 4970 4660 4990 4700
rect 5110 4660 5130 4700
rect 5250 4660 5270 4700
rect 5390 4660 5410 4700
rect 5530 4660 5550 4700
rect 5670 4660 5690 4700
rect 6020 5190 6040 5210
rect 6260 5190 6280 5210
rect 6610 5700 6630 5740
rect 6750 5700 6770 5740
rect 6890 5700 6910 5740
rect 7030 5700 7050 5740
rect 7170 5700 7190 5740
rect 7310 5700 7330 5740
rect 7450 5700 7470 5740
rect 7590 5700 7610 5740
rect 7730 5700 7750 5740
rect 7870 5700 7890 5740
rect 8010 5700 8030 5740
rect 5810 4660 5830 4700
rect 6020 4670 6040 4690
rect 6260 4670 6280 4690
rect 6470 4660 6490 4700
rect 6020 4190 6040 4210
rect 6260 4190 6280 4210
rect 6610 4660 6630 4700
rect 6750 4660 6770 4700
rect 6890 4660 6910 4700
rect 7030 4660 7050 4700
rect 7170 4660 7190 4700
rect 7310 4660 7330 4700
rect 7450 4660 7470 4700
rect 7590 4660 7610 4700
rect 7730 4660 7750 4700
rect 7870 4660 7890 4700
rect 8010 4660 8030 4700
rect 4240 3970 4280 3990
rect 4260 3430 4300 3450
rect 8020 3970 8060 3990
rect 8000 3430 8040 3450
rect 4260 2890 4300 2910
rect 8000 2890 8040 2910
<< psubdiff >>
rect 4460 7670 4490 7690
rect 4530 7670 4560 7690
rect 4460 7660 4560 7670
rect 4630 7670 4660 7690
rect 4700 7670 4730 7690
rect 4630 7660 4730 7670
rect 4800 7670 4830 7690
rect 4870 7670 4900 7690
rect 4800 7660 4900 7670
rect 4970 7670 5000 7690
rect 5040 7670 5070 7690
rect 4970 7660 5070 7670
rect 5140 7670 5170 7690
rect 5210 7670 5240 7690
rect 5140 7660 5240 7670
rect 5310 7670 5340 7690
rect 5380 7670 5410 7690
rect 5310 7660 5410 7670
rect 5480 7670 5510 7690
rect 5550 7670 5580 7690
rect 5480 7660 5580 7670
rect 5650 7670 5680 7690
rect 5720 7670 5750 7690
rect 5650 7660 5750 7670
rect 5820 7670 5850 7690
rect 5890 7670 5920 7690
rect 5820 7660 5920 7670
rect 5990 7670 6020 7690
rect 6060 7670 6090 7690
rect 5990 7660 6090 7670
rect 6210 7670 6240 7690
rect 6280 7670 6310 7690
rect 6210 7660 6310 7670
rect 6380 7670 6410 7690
rect 6450 7670 6480 7690
rect 6380 7660 6480 7670
rect 6550 7670 6580 7690
rect 6620 7670 6650 7690
rect 6550 7660 6650 7670
rect 6720 7670 6750 7690
rect 6790 7670 6820 7690
rect 6720 7660 6820 7670
rect 6890 7670 6920 7690
rect 6960 7670 6990 7690
rect 6890 7660 6990 7670
rect 7060 7670 7090 7690
rect 7130 7670 7160 7690
rect 7060 7660 7160 7670
rect 7230 7670 7260 7690
rect 7300 7670 7330 7690
rect 7230 7660 7330 7670
rect 7400 7670 7430 7690
rect 7470 7670 7500 7690
rect 7400 7660 7500 7670
rect 7570 7670 7600 7690
rect 7640 7670 7670 7690
rect 7570 7660 7670 7670
rect 7740 7670 7770 7690
rect 7810 7670 7840 7690
rect 7740 7660 7840 7670
rect 4460 2730 4560 2740
rect 4460 2710 4490 2730
rect 4530 2710 4560 2730
rect 4630 2730 4730 2740
rect 4630 2710 4660 2730
rect 4700 2710 4730 2730
rect 4800 2730 4900 2740
rect 4800 2710 4830 2730
rect 4870 2710 4900 2730
rect 4970 2730 5070 2740
rect 4970 2710 5000 2730
rect 5040 2710 5070 2730
rect 5140 2730 5240 2740
rect 5140 2710 5170 2730
rect 5210 2710 5240 2730
rect 5310 2730 5410 2740
rect 5310 2710 5340 2730
rect 5380 2710 5410 2730
rect 5480 2730 5580 2740
rect 5480 2710 5510 2730
rect 5550 2710 5580 2730
rect 5650 2730 5750 2740
rect 5650 2710 5680 2730
rect 5720 2710 5750 2730
rect 5820 2730 5920 2740
rect 5820 2710 5850 2730
rect 5890 2710 5920 2730
rect 5990 2730 6090 2740
rect 5990 2710 6020 2730
rect 6060 2710 6090 2730
rect 6210 2730 6310 2740
rect 6210 2710 6240 2730
rect 6280 2710 6310 2730
rect 6380 2730 6480 2740
rect 6380 2710 6410 2730
rect 6450 2710 6480 2730
rect 6550 2730 6650 2740
rect 6550 2710 6580 2730
rect 6620 2710 6650 2730
rect 6720 2730 6820 2740
rect 6720 2710 6750 2730
rect 6790 2710 6820 2730
rect 6890 2730 6990 2740
rect 6890 2710 6920 2730
rect 6960 2710 6990 2730
rect 7060 2730 7160 2740
rect 7060 2710 7090 2730
rect 7130 2710 7160 2730
rect 7230 2730 7330 2740
rect 7230 2710 7260 2730
rect 7300 2710 7330 2730
rect 7400 2730 7500 2740
rect 7400 2710 7430 2730
rect 7470 2710 7500 2730
rect 7570 2730 7670 2740
rect 7570 2710 7600 2730
rect 7640 2710 7670 2730
rect 7740 2730 7840 2740
rect 7740 2710 7770 2730
rect 7810 2710 7840 2730
<< nsubdiff >>
rect 4220 6190 4260 6200
rect 4220 6150 4230 6190
rect 4250 6150 4260 6190
rect 4220 6140 4260 6150
rect 5900 5210 5960 5230
rect 5900 5190 5920 5210
rect 5940 5190 5960 5210
rect 4220 4250 4260 4260
rect 4220 4210 4230 4250
rect 4250 4210 4260 4250
rect 4220 4200 4260 4210
rect 5900 5170 5960 5190
rect 6340 5210 6400 5230
rect 8040 6190 8080 6200
rect 8040 6150 8050 6190
rect 8070 6150 8080 6190
rect 8040 6140 8080 6150
rect 6340 5190 6360 5210
rect 6380 5190 6400 5210
rect 6340 5170 6400 5190
rect 8040 4250 8080 4260
rect 8040 4210 8050 4250
rect 8070 4210 8080 4250
rect 8040 4200 8080 4210
<< psubdiffcont >>
rect 4490 7670 4530 7690
rect 4660 7670 4700 7690
rect 4830 7670 4870 7690
rect 5000 7670 5040 7690
rect 5170 7670 5210 7690
rect 5340 7670 5380 7690
rect 5510 7670 5550 7690
rect 5680 7670 5720 7690
rect 5850 7670 5890 7690
rect 6020 7670 6060 7690
rect 6240 7670 6280 7690
rect 6410 7670 6450 7690
rect 6580 7670 6620 7690
rect 6750 7670 6790 7690
rect 6920 7670 6960 7690
rect 7090 7670 7130 7690
rect 7260 7670 7300 7690
rect 7430 7670 7470 7690
rect 7600 7670 7640 7690
rect 7770 7670 7810 7690
rect 4490 2710 4530 2730
rect 4660 2710 4700 2730
rect 4830 2710 4870 2730
rect 5000 2710 5040 2730
rect 5170 2710 5210 2730
rect 5340 2710 5380 2730
rect 5510 2710 5550 2730
rect 5680 2710 5720 2730
rect 5850 2710 5890 2730
rect 6020 2710 6060 2730
rect 6240 2710 6280 2730
rect 6410 2710 6450 2730
rect 6580 2710 6620 2730
rect 6750 2710 6790 2730
rect 6920 2710 6960 2730
rect 7090 2710 7130 2730
rect 7260 2710 7300 2730
rect 7430 2710 7470 2730
rect 7600 2710 7640 2730
rect 7770 2710 7810 2730
<< nsubdiffcont >>
rect 4230 6150 4250 6190
rect 5920 5190 5940 5210
rect 4230 4210 4250 4250
rect 8050 6150 8070 6190
rect 6360 5190 6380 5210
rect 8050 4210 8070 4250
<< poly >>
rect 4400 7670 4440 7680
rect 4400 7650 4410 7670
rect 4430 7650 4440 7670
rect 4400 7620 4440 7650
rect 7860 7670 7900 7680
rect 7860 7650 7870 7670
rect 7890 7650 7900 7670
rect 7860 7620 7900 7650
rect 4150 7570 4190 7580
rect 4150 7550 4160 7570
rect 4180 7550 4190 7570
rect 4150 7540 4190 7550
rect 4150 7480 4170 7540
rect 4400 7520 4460 7620
rect 4560 7590 4580 7620
rect 4610 7590 4630 7620
rect 4560 7550 4630 7590
rect 4560 7520 4580 7550
rect 4610 7520 4630 7550
rect 4730 7590 4750 7620
rect 4780 7590 4800 7620
rect 4730 7550 4800 7590
rect 4730 7520 4750 7550
rect 4780 7520 4800 7550
rect 4900 7590 4920 7620
rect 4950 7590 4970 7620
rect 4900 7550 4970 7590
rect 4900 7520 4920 7550
rect 4950 7520 4970 7550
rect 5070 7590 5090 7620
rect 5120 7590 5140 7620
rect 5070 7550 5140 7590
rect 5070 7520 5090 7550
rect 5120 7520 5140 7550
rect 5240 7590 5260 7620
rect 5290 7590 5310 7620
rect 5240 7550 5310 7590
rect 5240 7520 5260 7550
rect 5290 7520 5310 7550
rect 5410 7590 5430 7620
rect 5460 7590 5480 7620
rect 5410 7550 5480 7590
rect 5410 7520 5430 7550
rect 5460 7520 5480 7550
rect 5580 7590 5600 7620
rect 5630 7590 5650 7620
rect 5580 7550 5650 7590
rect 5580 7520 5600 7550
rect 5630 7520 5650 7550
rect 5750 7590 5770 7620
rect 5800 7590 5820 7620
rect 5750 7550 5820 7590
rect 5750 7520 5770 7550
rect 5800 7520 5820 7550
rect 5920 7590 5940 7620
rect 5970 7590 5990 7620
rect 5920 7550 5990 7590
rect 5920 7520 5940 7550
rect 5970 7520 5990 7550
rect 6090 7590 6110 7620
rect 6190 7590 6210 7620
rect 6090 7550 6210 7590
rect 6090 7520 6110 7550
rect 6190 7520 6210 7550
rect 6310 7590 6330 7620
rect 6360 7590 6380 7620
rect 6310 7550 6380 7590
rect 6310 7520 6330 7550
rect 6360 7520 6380 7550
rect 6480 7590 6500 7620
rect 6530 7590 6550 7620
rect 6480 7550 6550 7590
rect 6480 7520 6500 7550
rect 6530 7520 6550 7550
rect 6650 7590 6670 7620
rect 6700 7590 6720 7620
rect 6650 7550 6720 7590
rect 6650 7520 6670 7550
rect 6700 7520 6720 7550
rect 6820 7590 6840 7620
rect 6870 7590 6890 7620
rect 6820 7550 6890 7590
rect 6820 7520 6840 7550
rect 6870 7520 6890 7550
rect 6990 7590 7010 7620
rect 7040 7590 7060 7620
rect 6990 7550 7060 7590
rect 6990 7520 7010 7550
rect 7040 7520 7060 7550
rect 7160 7590 7180 7620
rect 7210 7590 7230 7620
rect 7160 7550 7230 7590
rect 7160 7520 7180 7550
rect 7210 7520 7230 7550
rect 7330 7590 7350 7620
rect 7380 7590 7400 7620
rect 7330 7550 7400 7590
rect 7330 7520 7350 7550
rect 7380 7520 7400 7550
rect 7500 7590 7520 7620
rect 7550 7590 7570 7620
rect 7500 7550 7570 7590
rect 7500 7520 7520 7550
rect 7550 7520 7570 7550
rect 7670 7590 7690 7620
rect 7720 7590 7740 7620
rect 7670 7550 7740 7590
rect 7670 7520 7690 7550
rect 7720 7520 7740 7550
rect 7840 7520 7900 7620
rect 8110 7570 8150 7580
rect 8110 7550 8120 7570
rect 8140 7550 8150 7570
rect 8110 7540 8150 7550
rect 8130 7480 8150 7540
rect 4150 6980 4180 7480
rect 4380 6980 4400 7480
rect 4440 7380 4460 7480
rect 4560 7450 4580 7480
rect 4610 7450 4630 7480
rect 4560 7410 4630 7450
rect 4560 7380 4580 7410
rect 4610 7380 4630 7410
rect 4730 7450 4750 7480
rect 4780 7450 4800 7480
rect 4730 7410 4800 7450
rect 4730 7380 4750 7410
rect 4780 7380 4800 7410
rect 4900 7450 4920 7480
rect 4950 7450 4970 7480
rect 4900 7410 4970 7450
rect 4900 7380 4920 7410
rect 4950 7380 4970 7410
rect 5070 7450 5090 7480
rect 5120 7450 5140 7480
rect 5070 7410 5140 7450
rect 5070 7380 5090 7410
rect 5120 7380 5140 7410
rect 5240 7450 5260 7480
rect 5290 7450 5310 7480
rect 5240 7410 5310 7450
rect 5240 7380 5260 7410
rect 5290 7380 5310 7410
rect 5410 7450 5430 7480
rect 5460 7450 5480 7480
rect 5410 7410 5480 7450
rect 5410 7380 5430 7410
rect 5460 7380 5480 7410
rect 5580 7450 5600 7480
rect 5630 7450 5650 7480
rect 5580 7410 5650 7450
rect 5580 7380 5600 7410
rect 5630 7380 5650 7410
rect 5750 7450 5770 7480
rect 5800 7450 5820 7480
rect 5750 7410 5820 7450
rect 5750 7380 5770 7410
rect 5800 7380 5820 7410
rect 5920 7450 5940 7480
rect 5970 7450 5990 7480
rect 5920 7410 5990 7450
rect 5920 7380 5940 7410
rect 5970 7380 5990 7410
rect 6090 7450 6110 7480
rect 6190 7450 6210 7480
rect 6090 7410 6210 7450
rect 6090 7380 6110 7410
rect 4160 6440 4180 6940
rect 4380 6440 4410 6940
rect 4390 6380 4410 6440
rect 4370 6370 4410 6380
rect 4370 6350 4380 6370
rect 4400 6350 4410 6370
rect 4370 6340 4410 6350
rect 4440 6340 4460 7340
rect 4560 7310 4580 7340
rect 4610 7310 4630 7340
rect 4560 7270 4630 7310
rect 4560 7210 4580 7270
rect 4610 7210 4630 7270
rect 4560 7170 4630 7210
rect 4560 7110 4580 7170
rect 4610 7110 4630 7170
rect 4560 7070 4630 7110
rect 4560 7010 4580 7070
rect 4610 7010 4630 7070
rect 4560 6970 4630 7010
rect 4560 6910 4580 6970
rect 4610 6910 4630 6970
rect 4560 6870 4630 6910
rect 4560 6810 4580 6870
rect 4610 6810 4630 6870
rect 4560 6770 4630 6810
rect 4560 6710 4580 6770
rect 4610 6710 4630 6770
rect 4560 6670 4630 6710
rect 4560 6610 4580 6670
rect 4610 6610 4630 6670
rect 4560 6570 4630 6610
rect 4560 6510 4580 6570
rect 4610 6510 4630 6570
rect 4560 6470 4630 6510
rect 4560 6410 4580 6470
rect 4610 6410 4630 6470
rect 4560 6370 4630 6410
rect 4560 6340 4580 6370
rect 4610 6340 4630 6370
rect 4730 7310 4750 7340
rect 4780 7310 4800 7340
rect 4730 7270 4800 7310
rect 4730 7210 4750 7270
rect 4780 7210 4800 7270
rect 4730 7170 4800 7210
rect 4730 7110 4750 7170
rect 4780 7110 4800 7170
rect 4730 7070 4800 7110
rect 4730 7010 4750 7070
rect 4780 7010 4800 7070
rect 4730 6970 4800 7010
rect 4730 6910 4750 6970
rect 4780 6910 4800 6970
rect 4730 6870 4800 6910
rect 4730 6810 4750 6870
rect 4780 6810 4800 6870
rect 4730 6770 4800 6810
rect 4730 6710 4750 6770
rect 4780 6710 4800 6770
rect 4730 6670 4800 6710
rect 4730 6610 4750 6670
rect 4780 6610 4800 6670
rect 4730 6570 4800 6610
rect 4730 6510 4750 6570
rect 4780 6510 4800 6570
rect 4730 6470 4800 6510
rect 4730 6410 4750 6470
rect 4780 6410 4800 6470
rect 4730 6370 4800 6410
rect 4730 6340 4750 6370
rect 4780 6340 4800 6370
rect 4900 7310 4920 7340
rect 4950 7310 4970 7340
rect 4900 7270 4970 7310
rect 4900 7210 4920 7270
rect 4950 7210 4970 7270
rect 4900 7170 4970 7210
rect 4900 7110 4920 7170
rect 4950 7110 4970 7170
rect 4900 7070 4970 7110
rect 4900 7010 4920 7070
rect 4950 7010 4970 7070
rect 4900 6970 4970 7010
rect 4900 6910 4920 6970
rect 4950 6910 4970 6970
rect 4900 6870 4970 6910
rect 4900 6810 4920 6870
rect 4950 6810 4970 6870
rect 4900 6770 4970 6810
rect 4900 6710 4920 6770
rect 4950 6710 4970 6770
rect 4900 6670 4970 6710
rect 4900 6610 4920 6670
rect 4950 6610 4970 6670
rect 4900 6570 4970 6610
rect 4900 6510 4920 6570
rect 4950 6510 4970 6570
rect 4900 6470 4970 6510
rect 4900 6410 4920 6470
rect 4950 6410 4970 6470
rect 4900 6370 4970 6410
rect 4900 6340 4920 6370
rect 4950 6340 4970 6370
rect 5070 7310 5090 7340
rect 5120 7310 5140 7340
rect 5070 7270 5140 7310
rect 5070 7210 5090 7270
rect 5120 7210 5140 7270
rect 5070 7170 5140 7210
rect 5070 7110 5090 7170
rect 5120 7110 5140 7170
rect 5070 7070 5140 7110
rect 5070 7010 5090 7070
rect 5120 7010 5140 7070
rect 5070 6970 5140 7010
rect 5070 6910 5090 6970
rect 5120 6910 5140 6970
rect 5070 6870 5140 6910
rect 5070 6810 5090 6870
rect 5120 6810 5140 6870
rect 5070 6770 5140 6810
rect 5070 6710 5090 6770
rect 5120 6710 5140 6770
rect 5070 6670 5140 6710
rect 5070 6610 5090 6670
rect 5120 6610 5140 6670
rect 5070 6570 5140 6610
rect 5070 6510 5090 6570
rect 5120 6510 5140 6570
rect 5070 6470 5140 6510
rect 5070 6410 5090 6470
rect 5120 6410 5140 6470
rect 5070 6370 5140 6410
rect 5070 6340 5090 6370
rect 5120 6340 5140 6370
rect 5240 7310 5260 7340
rect 5290 7310 5310 7340
rect 5240 7270 5310 7310
rect 5240 7210 5260 7270
rect 5290 7210 5310 7270
rect 5240 7170 5310 7210
rect 5240 7110 5260 7170
rect 5290 7110 5310 7170
rect 5240 7070 5310 7110
rect 5240 7010 5260 7070
rect 5290 7010 5310 7070
rect 5240 6970 5310 7010
rect 5240 6910 5260 6970
rect 5290 6910 5310 6970
rect 5240 6870 5310 6910
rect 5240 6810 5260 6870
rect 5290 6810 5310 6870
rect 5240 6770 5310 6810
rect 5240 6710 5260 6770
rect 5290 6710 5310 6770
rect 5240 6670 5310 6710
rect 5240 6610 5260 6670
rect 5290 6610 5310 6670
rect 5240 6570 5310 6610
rect 5240 6510 5260 6570
rect 5290 6510 5310 6570
rect 5240 6470 5310 6510
rect 5240 6410 5260 6470
rect 5290 6410 5310 6470
rect 5240 6370 5310 6410
rect 5240 6340 5260 6370
rect 5290 6340 5310 6370
rect 5410 7310 5430 7340
rect 5460 7310 5480 7340
rect 5410 7270 5480 7310
rect 5410 7210 5430 7270
rect 5460 7210 5480 7270
rect 5410 7170 5480 7210
rect 5410 7110 5430 7170
rect 5460 7110 5480 7170
rect 5410 7070 5480 7110
rect 5410 7010 5430 7070
rect 5460 7010 5480 7070
rect 5410 6970 5480 7010
rect 5410 6910 5430 6970
rect 5460 6910 5480 6970
rect 5410 6870 5480 6910
rect 5410 6810 5430 6870
rect 5460 6810 5480 6870
rect 5410 6770 5480 6810
rect 5410 6710 5430 6770
rect 5460 6710 5480 6770
rect 5410 6670 5480 6710
rect 5410 6610 5430 6670
rect 5460 6610 5480 6670
rect 5410 6570 5480 6610
rect 5410 6510 5430 6570
rect 5460 6510 5480 6570
rect 5410 6470 5480 6510
rect 5410 6410 5430 6470
rect 5460 6410 5480 6470
rect 5410 6370 5480 6410
rect 5410 6340 5430 6370
rect 5460 6340 5480 6370
rect 5580 7310 5600 7340
rect 5630 7310 5650 7340
rect 5580 7270 5650 7310
rect 5580 7210 5600 7270
rect 5630 7210 5650 7270
rect 5580 7170 5650 7210
rect 5580 7110 5600 7170
rect 5630 7110 5650 7170
rect 5580 7070 5650 7110
rect 5580 7010 5600 7070
rect 5630 7010 5650 7070
rect 5580 6970 5650 7010
rect 5580 6910 5600 6970
rect 5630 6910 5650 6970
rect 5580 6870 5650 6910
rect 5580 6810 5600 6870
rect 5630 6810 5650 6870
rect 5580 6770 5650 6810
rect 5580 6710 5600 6770
rect 5630 6710 5650 6770
rect 5580 6670 5650 6710
rect 5580 6610 5600 6670
rect 5630 6610 5650 6670
rect 5580 6570 5650 6610
rect 5580 6510 5600 6570
rect 5630 6510 5650 6570
rect 5580 6470 5650 6510
rect 5580 6410 5600 6470
rect 5630 6410 5650 6470
rect 5580 6370 5650 6410
rect 5580 6340 5600 6370
rect 5630 6340 5650 6370
rect 5750 7310 5770 7340
rect 5800 7310 5820 7340
rect 5750 7270 5820 7310
rect 5750 7210 5770 7270
rect 5800 7210 5820 7270
rect 5750 7170 5820 7210
rect 5750 7110 5770 7170
rect 5800 7110 5820 7170
rect 5750 7070 5820 7110
rect 5750 7010 5770 7070
rect 5800 7010 5820 7070
rect 5750 6970 5820 7010
rect 5750 6910 5770 6970
rect 5800 6910 5820 6970
rect 5750 6870 5820 6910
rect 5750 6810 5770 6870
rect 5800 6810 5820 6870
rect 5750 6770 5820 6810
rect 5750 6710 5770 6770
rect 5800 6710 5820 6770
rect 5750 6670 5820 6710
rect 5750 6610 5770 6670
rect 5800 6610 5820 6670
rect 5750 6570 5820 6610
rect 5750 6510 5770 6570
rect 5800 6510 5820 6570
rect 5750 6470 5820 6510
rect 5750 6410 5770 6470
rect 5800 6410 5820 6470
rect 5750 6370 5820 6410
rect 5750 6340 5770 6370
rect 5800 6340 5820 6370
rect 5920 7310 5940 7340
rect 5970 7310 5990 7340
rect 5920 7270 5990 7310
rect 5920 7210 5940 7270
rect 5970 7210 5990 7270
rect 5920 7170 5990 7210
rect 5920 7110 5940 7170
rect 5970 7110 5990 7170
rect 5920 7070 5990 7110
rect 5920 7010 5940 7070
rect 5970 7010 5990 7070
rect 5920 6970 5990 7010
rect 5920 6910 5940 6970
rect 5970 6910 5990 6970
rect 5920 6870 5990 6910
rect 5920 6810 5940 6870
rect 5970 6810 5990 6870
rect 5920 6770 5990 6810
rect 5920 6710 5940 6770
rect 5970 6710 5990 6770
rect 5920 6670 5990 6710
rect 5920 6610 5940 6670
rect 5970 6610 5990 6670
rect 5920 6570 5990 6610
rect 5920 6510 5940 6570
rect 5970 6510 5990 6570
rect 5920 6470 5990 6510
rect 5920 6410 5940 6470
rect 5970 6410 5990 6470
rect 5920 6370 5990 6410
rect 5920 6340 5940 6370
rect 5970 6340 5990 6370
rect 6090 7310 6110 7340
rect 6140 7310 6160 7410
rect 6190 7380 6210 7410
rect 6310 7450 6330 7480
rect 6360 7450 6380 7480
rect 6310 7410 6380 7450
rect 6310 7380 6330 7410
rect 6360 7380 6380 7410
rect 6480 7450 6500 7480
rect 6530 7450 6550 7480
rect 6480 7410 6550 7450
rect 6480 7380 6500 7410
rect 6530 7380 6550 7410
rect 6650 7450 6670 7480
rect 6700 7450 6720 7480
rect 6650 7410 6720 7450
rect 6650 7380 6670 7410
rect 6700 7380 6720 7410
rect 6820 7450 6840 7480
rect 6870 7450 6890 7480
rect 6820 7410 6890 7450
rect 6820 7380 6840 7410
rect 6870 7380 6890 7410
rect 6990 7450 7010 7480
rect 7040 7450 7060 7480
rect 6990 7410 7060 7450
rect 6990 7380 7010 7410
rect 7040 7380 7060 7410
rect 7160 7450 7180 7480
rect 7210 7450 7230 7480
rect 7160 7410 7230 7450
rect 7160 7380 7180 7410
rect 7210 7380 7230 7410
rect 7330 7450 7350 7480
rect 7380 7450 7400 7480
rect 7330 7410 7400 7450
rect 7330 7380 7350 7410
rect 7380 7380 7400 7410
rect 7500 7450 7520 7480
rect 7550 7450 7570 7480
rect 7500 7410 7570 7450
rect 7500 7380 7520 7410
rect 7550 7380 7570 7410
rect 7670 7450 7690 7480
rect 7720 7450 7740 7480
rect 7670 7410 7740 7450
rect 7670 7380 7690 7410
rect 7720 7380 7740 7410
rect 7840 7380 7860 7480
rect 6190 7310 6210 7340
rect 6090 7270 6210 7310
rect 6090 7210 6110 7270
rect 6140 7210 6160 7270
rect 6190 7210 6210 7270
rect 6090 7170 6210 7210
rect 6090 7110 6110 7170
rect 6140 7110 6160 7170
rect 6190 7110 6210 7170
rect 6090 7070 6210 7110
rect 6090 7010 6110 7070
rect 6140 7010 6160 7070
rect 6190 7010 6210 7070
rect 6090 6970 6210 7010
rect 6090 6910 6110 6970
rect 6140 6910 6160 6970
rect 6190 6910 6210 6970
rect 6090 6870 6210 6910
rect 6090 6810 6110 6870
rect 6140 6810 6160 6870
rect 6190 6810 6210 6870
rect 6090 6770 6210 6810
rect 6090 6710 6110 6770
rect 6140 6710 6160 6770
rect 6190 6710 6210 6770
rect 6090 6670 6210 6710
rect 6090 6610 6110 6670
rect 6140 6610 6160 6670
rect 6190 6610 6210 6670
rect 6090 6570 6210 6610
rect 6090 6510 6110 6570
rect 6140 6510 6160 6570
rect 6190 6510 6210 6570
rect 6090 6470 6210 6510
rect 6090 6410 6110 6470
rect 6140 6410 6160 6470
rect 6190 6410 6210 6470
rect 6090 6370 6210 6410
rect 6090 6340 6110 6370
rect 6140 6280 6160 6370
rect 6190 6340 6210 6370
rect 6310 7310 6330 7340
rect 6360 7310 6380 7340
rect 6310 7270 6380 7310
rect 6310 7210 6330 7270
rect 6360 7210 6380 7270
rect 6310 7170 6380 7210
rect 6310 7110 6330 7170
rect 6360 7110 6380 7170
rect 6310 7070 6380 7110
rect 6310 7010 6330 7070
rect 6360 7010 6380 7070
rect 6310 6970 6380 7010
rect 6310 6910 6330 6970
rect 6360 6910 6380 6970
rect 6310 6870 6380 6910
rect 6310 6810 6330 6870
rect 6360 6810 6380 6870
rect 6310 6770 6380 6810
rect 6310 6710 6330 6770
rect 6360 6710 6380 6770
rect 6310 6670 6380 6710
rect 6310 6610 6330 6670
rect 6360 6610 6380 6670
rect 6310 6570 6380 6610
rect 6310 6510 6330 6570
rect 6360 6510 6380 6570
rect 6310 6470 6380 6510
rect 6310 6410 6330 6470
rect 6360 6410 6380 6470
rect 6310 6370 6380 6410
rect 6310 6340 6330 6370
rect 6360 6340 6380 6370
rect 6480 7310 6500 7340
rect 6530 7310 6550 7340
rect 6480 7270 6550 7310
rect 6480 7210 6500 7270
rect 6530 7210 6550 7270
rect 6480 7170 6550 7210
rect 6480 7110 6500 7170
rect 6530 7110 6550 7170
rect 6480 7070 6550 7110
rect 6480 7010 6500 7070
rect 6530 7010 6550 7070
rect 6480 6970 6550 7010
rect 6480 6910 6500 6970
rect 6530 6910 6550 6970
rect 6480 6870 6550 6910
rect 6480 6810 6500 6870
rect 6530 6810 6550 6870
rect 6480 6770 6550 6810
rect 6480 6710 6500 6770
rect 6530 6710 6550 6770
rect 6480 6670 6550 6710
rect 6480 6610 6500 6670
rect 6530 6610 6550 6670
rect 6480 6570 6550 6610
rect 6480 6510 6500 6570
rect 6530 6510 6550 6570
rect 6480 6470 6550 6510
rect 6480 6410 6500 6470
rect 6530 6410 6550 6470
rect 6480 6370 6550 6410
rect 6480 6340 6500 6370
rect 6530 6340 6550 6370
rect 6650 7310 6670 7340
rect 6700 7310 6720 7340
rect 6650 7270 6720 7310
rect 6650 7210 6670 7270
rect 6700 7210 6720 7270
rect 6650 7170 6720 7210
rect 6650 7110 6670 7170
rect 6700 7110 6720 7170
rect 6650 7070 6720 7110
rect 6650 7010 6670 7070
rect 6700 7010 6720 7070
rect 6650 6970 6720 7010
rect 6650 6910 6670 6970
rect 6700 6910 6720 6970
rect 6650 6870 6720 6910
rect 6650 6810 6670 6870
rect 6700 6810 6720 6870
rect 6650 6770 6720 6810
rect 6650 6710 6670 6770
rect 6700 6710 6720 6770
rect 6650 6670 6720 6710
rect 6650 6610 6670 6670
rect 6700 6610 6720 6670
rect 6650 6570 6720 6610
rect 6650 6510 6670 6570
rect 6700 6510 6720 6570
rect 6650 6470 6720 6510
rect 6650 6410 6670 6470
rect 6700 6410 6720 6470
rect 6650 6370 6720 6410
rect 6650 6340 6670 6370
rect 6700 6340 6720 6370
rect 6820 7310 6840 7340
rect 6870 7310 6890 7340
rect 6820 7270 6890 7310
rect 6820 7210 6840 7270
rect 6870 7210 6890 7270
rect 6820 7170 6890 7210
rect 6820 7110 6840 7170
rect 6870 7110 6890 7170
rect 6820 7070 6890 7110
rect 6820 7010 6840 7070
rect 6870 7010 6890 7070
rect 6820 6970 6890 7010
rect 6820 6910 6840 6970
rect 6870 6910 6890 6970
rect 6820 6870 6890 6910
rect 6820 6810 6840 6870
rect 6870 6810 6890 6870
rect 6820 6770 6890 6810
rect 6820 6710 6840 6770
rect 6870 6710 6890 6770
rect 6820 6670 6890 6710
rect 6820 6610 6840 6670
rect 6870 6610 6890 6670
rect 6820 6570 6890 6610
rect 6820 6510 6840 6570
rect 6870 6510 6890 6570
rect 6820 6470 6890 6510
rect 6820 6410 6840 6470
rect 6870 6410 6890 6470
rect 6820 6370 6890 6410
rect 6820 6340 6840 6370
rect 6870 6340 6890 6370
rect 6990 7310 7010 7340
rect 7040 7310 7060 7340
rect 6990 7270 7060 7310
rect 6990 7210 7010 7270
rect 7040 7210 7060 7270
rect 6990 7170 7060 7210
rect 6990 7110 7010 7170
rect 7040 7110 7060 7170
rect 6990 7070 7060 7110
rect 6990 7010 7010 7070
rect 7040 7010 7060 7070
rect 6990 6970 7060 7010
rect 6990 6910 7010 6970
rect 7040 6910 7060 6970
rect 6990 6870 7060 6910
rect 6990 6810 7010 6870
rect 7040 6810 7060 6870
rect 6990 6770 7060 6810
rect 6990 6710 7010 6770
rect 7040 6710 7060 6770
rect 6990 6670 7060 6710
rect 6990 6610 7010 6670
rect 7040 6610 7060 6670
rect 6990 6570 7060 6610
rect 6990 6510 7010 6570
rect 7040 6510 7060 6570
rect 6990 6470 7060 6510
rect 6990 6410 7010 6470
rect 7040 6410 7060 6470
rect 6990 6370 7060 6410
rect 6990 6340 7010 6370
rect 7040 6340 7060 6370
rect 7160 7310 7180 7340
rect 7210 7310 7230 7340
rect 7160 7270 7230 7310
rect 7160 7210 7180 7270
rect 7210 7210 7230 7270
rect 7160 7170 7230 7210
rect 7160 7110 7180 7170
rect 7210 7110 7230 7170
rect 7160 7070 7230 7110
rect 7160 7010 7180 7070
rect 7210 7010 7230 7070
rect 7160 6970 7230 7010
rect 7160 6910 7180 6970
rect 7210 6910 7230 6970
rect 7160 6870 7230 6910
rect 7160 6810 7180 6870
rect 7210 6810 7230 6870
rect 7160 6770 7230 6810
rect 7160 6710 7180 6770
rect 7210 6710 7230 6770
rect 7160 6670 7230 6710
rect 7160 6610 7180 6670
rect 7210 6610 7230 6670
rect 7160 6570 7230 6610
rect 7160 6510 7180 6570
rect 7210 6510 7230 6570
rect 7160 6470 7230 6510
rect 7160 6410 7180 6470
rect 7210 6410 7230 6470
rect 7160 6370 7230 6410
rect 7160 6340 7180 6370
rect 7210 6340 7230 6370
rect 7330 7310 7350 7340
rect 7380 7310 7400 7340
rect 7330 7270 7400 7310
rect 7330 7210 7350 7270
rect 7380 7210 7400 7270
rect 7330 7170 7400 7210
rect 7330 7110 7350 7170
rect 7380 7110 7400 7170
rect 7330 7070 7400 7110
rect 7330 7010 7350 7070
rect 7380 7010 7400 7070
rect 7330 6970 7400 7010
rect 7330 6910 7350 6970
rect 7380 6910 7400 6970
rect 7330 6870 7400 6910
rect 7330 6810 7350 6870
rect 7380 6810 7400 6870
rect 7330 6770 7400 6810
rect 7330 6710 7350 6770
rect 7380 6710 7400 6770
rect 7330 6670 7400 6710
rect 7330 6610 7350 6670
rect 7380 6610 7400 6670
rect 7330 6570 7400 6610
rect 7330 6510 7350 6570
rect 7380 6510 7400 6570
rect 7330 6470 7400 6510
rect 7330 6410 7350 6470
rect 7380 6410 7400 6470
rect 7330 6370 7400 6410
rect 7330 6340 7350 6370
rect 7380 6340 7400 6370
rect 7500 7310 7520 7340
rect 7550 7310 7570 7340
rect 7500 7270 7570 7310
rect 7500 7210 7520 7270
rect 7550 7210 7570 7270
rect 7500 7170 7570 7210
rect 7500 7110 7520 7170
rect 7550 7110 7570 7170
rect 7500 7070 7570 7110
rect 7500 7010 7520 7070
rect 7550 7010 7570 7070
rect 7500 6970 7570 7010
rect 7500 6910 7520 6970
rect 7550 6910 7570 6970
rect 7500 6870 7570 6910
rect 7500 6810 7520 6870
rect 7550 6810 7570 6870
rect 7500 6770 7570 6810
rect 7500 6710 7520 6770
rect 7550 6710 7570 6770
rect 7500 6670 7570 6710
rect 7500 6610 7520 6670
rect 7550 6610 7570 6670
rect 7500 6570 7570 6610
rect 7500 6510 7520 6570
rect 7550 6510 7570 6570
rect 7500 6470 7570 6510
rect 7500 6410 7520 6470
rect 7550 6410 7570 6470
rect 7500 6370 7570 6410
rect 7500 6340 7520 6370
rect 7550 6340 7570 6370
rect 7670 7310 7690 7340
rect 7720 7310 7740 7340
rect 7670 7270 7740 7310
rect 7670 7210 7690 7270
rect 7720 7210 7740 7270
rect 7670 7170 7740 7210
rect 7670 7110 7690 7170
rect 7720 7110 7740 7170
rect 7670 7070 7740 7110
rect 7670 7010 7690 7070
rect 7720 7010 7740 7070
rect 7670 6970 7740 7010
rect 7670 6910 7690 6970
rect 7720 6910 7740 6970
rect 7670 6870 7740 6910
rect 7670 6810 7690 6870
rect 7720 6810 7740 6870
rect 7670 6770 7740 6810
rect 7670 6710 7690 6770
rect 7720 6710 7740 6770
rect 7670 6670 7740 6710
rect 7670 6610 7690 6670
rect 7720 6610 7740 6670
rect 7670 6570 7740 6610
rect 7670 6510 7690 6570
rect 7720 6510 7740 6570
rect 7670 6470 7740 6510
rect 7670 6410 7690 6470
rect 7720 6410 7740 6470
rect 7670 6370 7740 6410
rect 7670 6340 7690 6370
rect 7720 6340 7740 6370
rect 7840 6340 7860 7340
rect 7900 6980 7920 7480
rect 8120 6980 8150 7480
rect 7890 6440 7920 6940
rect 8120 6440 8140 6940
rect 7890 6380 7910 6440
rect 7890 6370 7930 6380
rect 7890 6350 7900 6370
rect 7920 6350 7930 6370
rect 7890 6340 7930 6350
rect 4250 6270 4400 6280
rect 4250 6250 4260 6270
rect 4280 6250 4400 6270
rect 4250 6240 4400 6250
rect 4300 6220 4400 6240
rect 4440 6270 4680 6280
rect 4440 6250 4550 6270
rect 4570 6250 4680 6270
rect 4440 6240 4680 6250
rect 4440 6220 4540 6240
rect 4580 6220 4680 6240
rect 4720 6270 4960 6280
rect 4720 6250 4830 6270
rect 4850 6250 4960 6270
rect 4720 6240 4960 6250
rect 4720 6220 4820 6240
rect 4860 6220 4960 6240
rect 5000 6270 5240 6280
rect 5000 6250 5110 6270
rect 5130 6250 5240 6270
rect 5000 6240 5240 6250
rect 5000 6220 5100 6240
rect 5140 6220 5240 6240
rect 5280 6270 5520 6280
rect 5280 6250 5390 6270
rect 5410 6250 5520 6270
rect 5280 6240 5520 6250
rect 5280 6220 5380 6240
rect 5420 6220 5520 6240
rect 5560 6270 5800 6280
rect 5560 6250 5670 6270
rect 5690 6250 5800 6270
rect 5560 6240 5800 6250
rect 6070 6270 6230 6280
rect 6070 6250 6080 6270
rect 6100 6250 6200 6270
rect 6220 6250 6230 6270
rect 6070 6240 6230 6250
rect 6500 6270 6740 6280
rect 6500 6250 6610 6270
rect 6630 6250 6740 6270
rect 6500 6240 6740 6250
rect 5560 6220 5660 6240
rect 5700 6220 5800 6240
rect 6500 6220 6600 6240
rect 6640 6220 6740 6240
rect 6780 6270 7020 6280
rect 6780 6250 6890 6270
rect 6910 6250 7020 6270
rect 6780 6240 7020 6250
rect 6780 6220 6880 6240
rect 6920 6220 7020 6240
rect 7060 6270 7300 6280
rect 7060 6250 7170 6270
rect 7190 6250 7300 6270
rect 7060 6240 7300 6250
rect 7060 6220 7160 6240
rect 7200 6220 7300 6240
rect 7340 6270 7580 6280
rect 7340 6250 7450 6270
rect 7470 6250 7580 6270
rect 7340 6240 7580 6250
rect 7340 6220 7440 6240
rect 7480 6220 7580 6240
rect 7620 6270 7860 6280
rect 7620 6250 7730 6270
rect 7750 6250 7860 6270
rect 7620 6240 7860 6250
rect 7620 6220 7720 6240
rect 7760 6220 7860 6240
rect 7900 6270 8050 6280
rect 7900 6250 8020 6270
rect 8040 6250 8050 6270
rect 7900 6240 8050 6250
rect 7900 6220 8000 6240
rect 4300 5180 4400 5220
rect 4440 5180 4540 5220
rect 4580 5180 4680 5220
rect 4720 5180 4820 5220
rect 4860 5180 4960 5220
rect 5000 5180 5100 5220
rect 5140 5180 5240 5220
rect 5280 5180 5380 5220
rect 5420 5180 5520 5220
rect 5560 5180 5660 5220
rect 5700 5180 5800 5220
rect 6500 5180 6600 5220
rect 6640 5180 6740 5220
rect 6780 5180 6880 5220
rect 6920 5180 7020 5220
rect 7060 5180 7160 5220
rect 7200 5180 7300 5220
rect 7340 5180 7440 5220
rect 7480 5180 7580 5220
rect 7620 5180 7720 5220
rect 7760 5180 7860 5220
rect 7900 5180 8000 5220
rect 4300 4160 4400 4180
rect 4250 4150 4400 4160
rect 4250 4130 4260 4150
rect 4280 4130 4400 4150
rect 4250 4120 4400 4130
rect 4440 4160 4540 4180
rect 4580 4160 4680 4180
rect 4440 4150 4680 4160
rect 4440 4130 4550 4150
rect 4570 4130 4680 4150
rect 4440 4120 4680 4130
rect 4720 4160 4820 4180
rect 4860 4160 4960 4180
rect 4720 4150 4960 4160
rect 4720 4130 4830 4150
rect 4850 4130 4960 4150
rect 4720 4120 4960 4130
rect 5000 4160 5100 4180
rect 5140 4160 5240 4180
rect 5000 4150 5240 4160
rect 5000 4130 5110 4150
rect 5130 4130 5240 4150
rect 5000 4120 5240 4130
rect 5280 4160 5380 4180
rect 5420 4160 5520 4180
rect 5280 4150 5520 4160
rect 5280 4130 5390 4150
rect 5410 4130 5520 4150
rect 5280 4120 5520 4130
rect 5560 4160 5660 4180
rect 5700 4160 5800 4180
rect 6500 4160 6600 4180
rect 6640 4160 6740 4180
rect 5560 4150 5800 4160
rect 5560 4130 5670 4150
rect 5690 4130 5800 4150
rect 5560 4120 5800 4130
rect 6070 4150 6230 4160
rect 6070 4130 6080 4150
rect 6100 4130 6200 4150
rect 6220 4130 6230 4150
rect 6070 4120 6230 4130
rect 6500 4150 6740 4160
rect 6500 4130 6610 4150
rect 6630 4130 6740 4150
rect 6500 4120 6740 4130
rect 6780 4160 6880 4180
rect 6920 4160 7020 4180
rect 6780 4150 7020 4160
rect 6780 4130 6890 4150
rect 6910 4130 7020 4150
rect 6780 4120 7020 4130
rect 7060 4160 7160 4180
rect 7200 4160 7300 4180
rect 7060 4150 7300 4160
rect 7060 4130 7170 4150
rect 7190 4130 7300 4150
rect 7060 4120 7300 4130
rect 7340 4160 7440 4180
rect 7480 4160 7580 4180
rect 7340 4150 7580 4160
rect 7340 4130 7450 4150
rect 7470 4130 7580 4150
rect 7340 4120 7580 4130
rect 7620 4160 7720 4180
rect 7760 4160 7860 4180
rect 7620 4150 7860 4160
rect 7620 4130 7730 4150
rect 7750 4130 7860 4150
rect 7620 4120 7860 4130
rect 7900 4160 8000 4180
rect 7900 4150 8050 4160
rect 7900 4130 8020 4150
rect 8040 4130 8050 4150
rect 7900 4120 8050 4130
rect 4370 4050 4410 4060
rect 4370 4030 4380 4050
rect 4400 4030 4410 4050
rect 4370 4020 4410 4030
rect 4390 3960 4410 4020
rect 4160 3460 4180 3960
rect 4380 3460 4410 3960
rect 4150 2920 4180 3420
rect 4380 2920 4400 3420
rect 4440 3060 4460 4060
rect 4560 4030 4580 4060
rect 4610 4030 4630 4060
rect 4560 3990 4630 4030
rect 4560 3930 4580 3990
rect 4610 3930 4630 3990
rect 4560 3890 4630 3930
rect 4560 3830 4580 3890
rect 4610 3830 4630 3890
rect 4560 3790 4630 3830
rect 4560 3730 4580 3790
rect 4610 3730 4630 3790
rect 4560 3690 4630 3730
rect 4560 3630 4580 3690
rect 4610 3630 4630 3690
rect 4560 3590 4630 3630
rect 4560 3530 4580 3590
rect 4610 3530 4630 3590
rect 4560 3490 4630 3530
rect 4560 3430 4580 3490
rect 4610 3430 4630 3490
rect 4560 3390 4630 3430
rect 4560 3330 4580 3390
rect 4610 3330 4630 3390
rect 4560 3290 4630 3330
rect 4560 3230 4580 3290
rect 4610 3230 4630 3290
rect 4560 3190 4630 3230
rect 4560 3130 4580 3190
rect 4610 3130 4630 3190
rect 4560 3090 4630 3130
rect 4560 3060 4580 3090
rect 4610 3060 4630 3090
rect 4730 4030 4750 4060
rect 4780 4030 4800 4060
rect 4730 3990 4800 4030
rect 4730 3930 4750 3990
rect 4780 3930 4800 3990
rect 4730 3890 4800 3930
rect 4730 3830 4750 3890
rect 4780 3830 4800 3890
rect 4730 3790 4800 3830
rect 4730 3730 4750 3790
rect 4780 3730 4800 3790
rect 4730 3690 4800 3730
rect 4730 3630 4750 3690
rect 4780 3630 4800 3690
rect 4730 3590 4800 3630
rect 4730 3530 4750 3590
rect 4780 3530 4800 3590
rect 4730 3490 4800 3530
rect 4730 3430 4750 3490
rect 4780 3430 4800 3490
rect 4730 3390 4800 3430
rect 4730 3330 4750 3390
rect 4780 3330 4800 3390
rect 4730 3290 4800 3330
rect 4730 3230 4750 3290
rect 4780 3230 4800 3290
rect 4730 3190 4800 3230
rect 4730 3130 4750 3190
rect 4780 3130 4800 3190
rect 4730 3090 4800 3130
rect 4730 3060 4750 3090
rect 4780 3060 4800 3090
rect 4900 4030 4920 4060
rect 4950 4030 4970 4060
rect 4900 3990 4970 4030
rect 4900 3930 4920 3990
rect 4950 3930 4970 3990
rect 4900 3890 4970 3930
rect 4900 3830 4920 3890
rect 4950 3830 4970 3890
rect 4900 3790 4970 3830
rect 4900 3730 4920 3790
rect 4950 3730 4970 3790
rect 4900 3690 4970 3730
rect 4900 3630 4920 3690
rect 4950 3630 4970 3690
rect 4900 3590 4970 3630
rect 4900 3530 4920 3590
rect 4950 3530 4970 3590
rect 4900 3490 4970 3530
rect 4900 3430 4920 3490
rect 4950 3430 4970 3490
rect 4900 3390 4970 3430
rect 4900 3330 4920 3390
rect 4950 3330 4970 3390
rect 4900 3290 4970 3330
rect 4900 3230 4920 3290
rect 4950 3230 4970 3290
rect 4900 3190 4970 3230
rect 4900 3130 4920 3190
rect 4950 3130 4970 3190
rect 4900 3090 4970 3130
rect 4900 3060 4920 3090
rect 4950 3060 4970 3090
rect 5070 4030 5090 4060
rect 5120 4030 5140 4060
rect 5070 3990 5140 4030
rect 5070 3930 5090 3990
rect 5120 3930 5140 3990
rect 5070 3890 5140 3930
rect 5070 3830 5090 3890
rect 5120 3830 5140 3890
rect 5070 3790 5140 3830
rect 5070 3730 5090 3790
rect 5120 3730 5140 3790
rect 5070 3690 5140 3730
rect 5070 3630 5090 3690
rect 5120 3630 5140 3690
rect 5070 3590 5140 3630
rect 5070 3530 5090 3590
rect 5120 3530 5140 3590
rect 5070 3490 5140 3530
rect 5070 3430 5090 3490
rect 5120 3430 5140 3490
rect 5070 3390 5140 3430
rect 5070 3330 5090 3390
rect 5120 3330 5140 3390
rect 5070 3290 5140 3330
rect 5070 3230 5090 3290
rect 5120 3230 5140 3290
rect 5070 3190 5140 3230
rect 5070 3130 5090 3190
rect 5120 3130 5140 3190
rect 5070 3090 5140 3130
rect 5070 3060 5090 3090
rect 5120 3060 5140 3090
rect 5240 4030 5260 4060
rect 5290 4030 5310 4060
rect 5240 3990 5310 4030
rect 5240 3930 5260 3990
rect 5290 3930 5310 3990
rect 5240 3890 5310 3930
rect 5240 3830 5260 3890
rect 5290 3830 5310 3890
rect 5240 3790 5310 3830
rect 5240 3730 5260 3790
rect 5290 3730 5310 3790
rect 5240 3690 5310 3730
rect 5240 3630 5260 3690
rect 5290 3630 5310 3690
rect 5240 3590 5310 3630
rect 5240 3530 5260 3590
rect 5290 3530 5310 3590
rect 5240 3490 5310 3530
rect 5240 3430 5260 3490
rect 5290 3430 5310 3490
rect 5240 3390 5310 3430
rect 5240 3330 5260 3390
rect 5290 3330 5310 3390
rect 5240 3290 5310 3330
rect 5240 3230 5260 3290
rect 5290 3230 5310 3290
rect 5240 3190 5310 3230
rect 5240 3130 5260 3190
rect 5290 3130 5310 3190
rect 5240 3090 5310 3130
rect 5240 3060 5260 3090
rect 5290 3060 5310 3090
rect 5410 4030 5430 4060
rect 5460 4030 5480 4060
rect 5410 3990 5480 4030
rect 5410 3930 5430 3990
rect 5460 3930 5480 3990
rect 5410 3890 5480 3930
rect 5410 3830 5430 3890
rect 5460 3830 5480 3890
rect 5410 3790 5480 3830
rect 5410 3730 5430 3790
rect 5460 3730 5480 3790
rect 5410 3690 5480 3730
rect 5410 3630 5430 3690
rect 5460 3630 5480 3690
rect 5410 3590 5480 3630
rect 5410 3530 5430 3590
rect 5460 3530 5480 3590
rect 5410 3490 5480 3530
rect 5410 3430 5430 3490
rect 5460 3430 5480 3490
rect 5410 3390 5480 3430
rect 5410 3330 5430 3390
rect 5460 3330 5480 3390
rect 5410 3290 5480 3330
rect 5410 3230 5430 3290
rect 5460 3230 5480 3290
rect 5410 3190 5480 3230
rect 5410 3130 5430 3190
rect 5460 3130 5480 3190
rect 5410 3090 5480 3130
rect 5410 3060 5430 3090
rect 5460 3060 5480 3090
rect 5580 4030 5600 4060
rect 5630 4030 5650 4060
rect 5580 3990 5650 4030
rect 5580 3930 5600 3990
rect 5630 3930 5650 3990
rect 5580 3890 5650 3930
rect 5580 3830 5600 3890
rect 5630 3830 5650 3890
rect 5580 3790 5650 3830
rect 5580 3730 5600 3790
rect 5630 3730 5650 3790
rect 5580 3690 5650 3730
rect 5580 3630 5600 3690
rect 5630 3630 5650 3690
rect 5580 3590 5650 3630
rect 5580 3530 5600 3590
rect 5630 3530 5650 3590
rect 5580 3490 5650 3530
rect 5580 3430 5600 3490
rect 5630 3430 5650 3490
rect 5580 3390 5650 3430
rect 5580 3330 5600 3390
rect 5630 3330 5650 3390
rect 5580 3290 5650 3330
rect 5580 3230 5600 3290
rect 5630 3230 5650 3290
rect 5580 3190 5650 3230
rect 5580 3130 5600 3190
rect 5630 3130 5650 3190
rect 5580 3090 5650 3130
rect 5580 3060 5600 3090
rect 5630 3060 5650 3090
rect 5750 4030 5770 4060
rect 5800 4030 5820 4060
rect 5750 3990 5820 4030
rect 5750 3930 5770 3990
rect 5800 3930 5820 3990
rect 5750 3890 5820 3930
rect 5750 3830 5770 3890
rect 5800 3830 5820 3890
rect 5750 3790 5820 3830
rect 5750 3730 5770 3790
rect 5800 3730 5820 3790
rect 5750 3690 5820 3730
rect 5750 3630 5770 3690
rect 5800 3630 5820 3690
rect 5750 3590 5820 3630
rect 5750 3530 5770 3590
rect 5800 3530 5820 3590
rect 5750 3490 5820 3530
rect 5750 3430 5770 3490
rect 5800 3430 5820 3490
rect 5750 3390 5820 3430
rect 5750 3330 5770 3390
rect 5800 3330 5820 3390
rect 5750 3290 5820 3330
rect 5750 3230 5770 3290
rect 5800 3230 5820 3290
rect 5750 3190 5820 3230
rect 5750 3130 5770 3190
rect 5800 3130 5820 3190
rect 5750 3090 5820 3130
rect 5750 3060 5770 3090
rect 5800 3060 5820 3090
rect 5920 4030 5940 4060
rect 5970 4030 5990 4060
rect 5920 3990 5990 4030
rect 5920 3930 5940 3990
rect 5970 3930 5990 3990
rect 5920 3890 5990 3930
rect 5920 3830 5940 3890
rect 5970 3830 5990 3890
rect 5920 3790 5990 3830
rect 5920 3730 5940 3790
rect 5970 3730 5990 3790
rect 5920 3690 5990 3730
rect 5920 3630 5940 3690
rect 5970 3630 5990 3690
rect 5920 3590 5990 3630
rect 5920 3530 5940 3590
rect 5970 3530 5990 3590
rect 5920 3490 5990 3530
rect 5920 3430 5940 3490
rect 5970 3430 5990 3490
rect 5920 3390 5990 3430
rect 5920 3330 5940 3390
rect 5970 3330 5990 3390
rect 5920 3290 5990 3330
rect 5920 3230 5940 3290
rect 5970 3230 5990 3290
rect 5920 3190 5990 3230
rect 5920 3130 5940 3190
rect 5970 3130 5990 3190
rect 5920 3090 5990 3130
rect 5920 3060 5940 3090
rect 5970 3060 5990 3090
rect 6090 4030 6110 4060
rect 6140 4030 6160 4120
rect 6190 4030 6210 4060
rect 6090 3990 6210 4030
rect 6090 3930 6110 3990
rect 6140 3930 6160 3990
rect 6190 3930 6210 3990
rect 6090 3890 6210 3930
rect 6090 3830 6110 3890
rect 6140 3830 6160 3890
rect 6190 3830 6210 3890
rect 6090 3790 6210 3830
rect 6090 3730 6110 3790
rect 6140 3730 6160 3790
rect 6190 3730 6210 3790
rect 6090 3690 6210 3730
rect 6090 3630 6110 3690
rect 6140 3630 6160 3690
rect 6190 3630 6210 3690
rect 6090 3590 6210 3630
rect 6090 3530 6110 3590
rect 6140 3530 6160 3590
rect 6190 3530 6210 3590
rect 6090 3490 6210 3530
rect 6090 3430 6110 3490
rect 6140 3430 6160 3490
rect 6190 3430 6210 3490
rect 6090 3390 6210 3430
rect 6090 3330 6110 3390
rect 6140 3330 6160 3390
rect 6190 3330 6210 3390
rect 6090 3290 6210 3330
rect 6090 3230 6110 3290
rect 6140 3230 6160 3290
rect 6190 3230 6210 3290
rect 6090 3190 6210 3230
rect 6090 3130 6110 3190
rect 6140 3130 6160 3190
rect 6190 3130 6210 3190
rect 6090 3090 6210 3130
rect 6090 3060 6110 3090
rect 4440 2920 4460 3020
rect 4560 2990 4580 3020
rect 4610 2990 4630 3020
rect 4560 2950 4630 2990
rect 4560 2920 4580 2950
rect 4610 2920 4630 2950
rect 4730 2990 4750 3020
rect 4780 2990 4800 3020
rect 4730 2950 4800 2990
rect 4730 2920 4750 2950
rect 4780 2920 4800 2950
rect 4900 2990 4920 3020
rect 4950 2990 4970 3020
rect 4900 2950 4970 2990
rect 4900 2920 4920 2950
rect 4950 2920 4970 2950
rect 5070 2990 5090 3020
rect 5120 2990 5140 3020
rect 5070 2950 5140 2990
rect 5070 2920 5090 2950
rect 5120 2920 5140 2950
rect 5240 2990 5260 3020
rect 5290 2990 5310 3020
rect 5240 2950 5310 2990
rect 5240 2920 5260 2950
rect 5290 2920 5310 2950
rect 5410 2990 5430 3020
rect 5460 2990 5480 3020
rect 5410 2950 5480 2990
rect 5410 2920 5430 2950
rect 5460 2920 5480 2950
rect 5580 2990 5600 3020
rect 5630 2990 5650 3020
rect 5580 2950 5650 2990
rect 5580 2920 5600 2950
rect 5630 2920 5650 2950
rect 5750 2990 5770 3020
rect 5800 2990 5820 3020
rect 5750 2950 5820 2990
rect 5750 2920 5770 2950
rect 5800 2920 5820 2950
rect 5920 2990 5940 3020
rect 5970 2990 5990 3020
rect 5920 2950 5990 2990
rect 5920 2920 5940 2950
rect 5970 2920 5990 2950
rect 6090 2990 6110 3020
rect 6140 2990 6160 3090
rect 6190 3060 6210 3090
rect 6310 4030 6330 4060
rect 6360 4030 6380 4060
rect 6310 3990 6380 4030
rect 6310 3930 6330 3990
rect 6360 3930 6380 3990
rect 6310 3890 6380 3930
rect 6310 3830 6330 3890
rect 6360 3830 6380 3890
rect 6310 3790 6380 3830
rect 6310 3730 6330 3790
rect 6360 3730 6380 3790
rect 6310 3690 6380 3730
rect 6310 3630 6330 3690
rect 6360 3630 6380 3690
rect 6310 3590 6380 3630
rect 6310 3530 6330 3590
rect 6360 3530 6380 3590
rect 6310 3490 6380 3530
rect 6310 3430 6330 3490
rect 6360 3430 6380 3490
rect 6310 3390 6380 3430
rect 6310 3330 6330 3390
rect 6360 3330 6380 3390
rect 6310 3290 6380 3330
rect 6310 3230 6330 3290
rect 6360 3230 6380 3290
rect 6310 3190 6380 3230
rect 6310 3130 6330 3190
rect 6360 3130 6380 3190
rect 6310 3090 6380 3130
rect 6310 3060 6330 3090
rect 6360 3060 6380 3090
rect 6480 4030 6500 4060
rect 6530 4030 6550 4060
rect 6480 3990 6550 4030
rect 6480 3930 6500 3990
rect 6530 3930 6550 3990
rect 6480 3890 6550 3930
rect 6480 3830 6500 3890
rect 6530 3830 6550 3890
rect 6480 3790 6550 3830
rect 6480 3730 6500 3790
rect 6530 3730 6550 3790
rect 6480 3690 6550 3730
rect 6480 3630 6500 3690
rect 6530 3630 6550 3690
rect 6480 3590 6550 3630
rect 6480 3530 6500 3590
rect 6530 3530 6550 3590
rect 6480 3490 6550 3530
rect 6480 3430 6500 3490
rect 6530 3430 6550 3490
rect 6480 3390 6550 3430
rect 6480 3330 6500 3390
rect 6530 3330 6550 3390
rect 6480 3290 6550 3330
rect 6480 3230 6500 3290
rect 6530 3230 6550 3290
rect 6480 3190 6550 3230
rect 6480 3130 6500 3190
rect 6530 3130 6550 3190
rect 6480 3090 6550 3130
rect 6480 3060 6500 3090
rect 6530 3060 6550 3090
rect 6650 4030 6670 4060
rect 6700 4030 6720 4060
rect 6650 3990 6720 4030
rect 6650 3930 6670 3990
rect 6700 3930 6720 3990
rect 6650 3890 6720 3930
rect 6650 3830 6670 3890
rect 6700 3830 6720 3890
rect 6650 3790 6720 3830
rect 6650 3730 6670 3790
rect 6700 3730 6720 3790
rect 6650 3690 6720 3730
rect 6650 3630 6670 3690
rect 6700 3630 6720 3690
rect 6650 3590 6720 3630
rect 6650 3530 6670 3590
rect 6700 3530 6720 3590
rect 6650 3490 6720 3530
rect 6650 3430 6670 3490
rect 6700 3430 6720 3490
rect 6650 3390 6720 3430
rect 6650 3330 6670 3390
rect 6700 3330 6720 3390
rect 6650 3290 6720 3330
rect 6650 3230 6670 3290
rect 6700 3230 6720 3290
rect 6650 3190 6720 3230
rect 6650 3130 6670 3190
rect 6700 3130 6720 3190
rect 6650 3090 6720 3130
rect 6650 3060 6670 3090
rect 6700 3060 6720 3090
rect 6820 4030 6840 4060
rect 6870 4030 6890 4060
rect 6820 3990 6890 4030
rect 6820 3930 6840 3990
rect 6870 3930 6890 3990
rect 6820 3890 6890 3930
rect 6820 3830 6840 3890
rect 6870 3830 6890 3890
rect 6820 3790 6890 3830
rect 6820 3730 6840 3790
rect 6870 3730 6890 3790
rect 6820 3690 6890 3730
rect 6820 3630 6840 3690
rect 6870 3630 6890 3690
rect 6820 3590 6890 3630
rect 6820 3530 6840 3590
rect 6870 3530 6890 3590
rect 6820 3490 6890 3530
rect 6820 3430 6840 3490
rect 6870 3430 6890 3490
rect 6820 3390 6890 3430
rect 6820 3330 6840 3390
rect 6870 3330 6890 3390
rect 6820 3290 6890 3330
rect 6820 3230 6840 3290
rect 6870 3230 6890 3290
rect 6820 3190 6890 3230
rect 6820 3130 6840 3190
rect 6870 3130 6890 3190
rect 6820 3090 6890 3130
rect 6820 3060 6840 3090
rect 6870 3060 6890 3090
rect 6990 4030 7010 4060
rect 7040 4030 7060 4060
rect 6990 3990 7060 4030
rect 6990 3930 7010 3990
rect 7040 3930 7060 3990
rect 6990 3890 7060 3930
rect 6990 3830 7010 3890
rect 7040 3830 7060 3890
rect 6990 3790 7060 3830
rect 6990 3730 7010 3790
rect 7040 3730 7060 3790
rect 6990 3690 7060 3730
rect 6990 3630 7010 3690
rect 7040 3630 7060 3690
rect 6990 3590 7060 3630
rect 6990 3530 7010 3590
rect 7040 3530 7060 3590
rect 6990 3490 7060 3530
rect 6990 3430 7010 3490
rect 7040 3430 7060 3490
rect 6990 3390 7060 3430
rect 6990 3330 7010 3390
rect 7040 3330 7060 3390
rect 6990 3290 7060 3330
rect 6990 3230 7010 3290
rect 7040 3230 7060 3290
rect 6990 3190 7060 3230
rect 6990 3130 7010 3190
rect 7040 3130 7060 3190
rect 6990 3090 7060 3130
rect 6990 3060 7010 3090
rect 7040 3060 7060 3090
rect 7160 4030 7180 4060
rect 7210 4030 7230 4060
rect 7160 3990 7230 4030
rect 7160 3930 7180 3990
rect 7210 3930 7230 3990
rect 7160 3890 7230 3930
rect 7160 3830 7180 3890
rect 7210 3830 7230 3890
rect 7160 3790 7230 3830
rect 7160 3730 7180 3790
rect 7210 3730 7230 3790
rect 7160 3690 7230 3730
rect 7160 3630 7180 3690
rect 7210 3630 7230 3690
rect 7160 3590 7230 3630
rect 7160 3530 7180 3590
rect 7210 3530 7230 3590
rect 7160 3490 7230 3530
rect 7160 3430 7180 3490
rect 7210 3430 7230 3490
rect 7160 3390 7230 3430
rect 7160 3330 7180 3390
rect 7210 3330 7230 3390
rect 7160 3290 7230 3330
rect 7160 3230 7180 3290
rect 7210 3230 7230 3290
rect 7160 3190 7230 3230
rect 7160 3130 7180 3190
rect 7210 3130 7230 3190
rect 7160 3090 7230 3130
rect 7160 3060 7180 3090
rect 7210 3060 7230 3090
rect 7330 4030 7350 4060
rect 7380 4030 7400 4060
rect 7330 3990 7400 4030
rect 7330 3930 7350 3990
rect 7380 3930 7400 3990
rect 7330 3890 7400 3930
rect 7330 3830 7350 3890
rect 7380 3830 7400 3890
rect 7330 3790 7400 3830
rect 7330 3730 7350 3790
rect 7380 3730 7400 3790
rect 7330 3690 7400 3730
rect 7330 3630 7350 3690
rect 7380 3630 7400 3690
rect 7330 3590 7400 3630
rect 7330 3530 7350 3590
rect 7380 3530 7400 3590
rect 7330 3490 7400 3530
rect 7330 3430 7350 3490
rect 7380 3430 7400 3490
rect 7330 3390 7400 3430
rect 7330 3330 7350 3390
rect 7380 3330 7400 3390
rect 7330 3290 7400 3330
rect 7330 3230 7350 3290
rect 7380 3230 7400 3290
rect 7330 3190 7400 3230
rect 7330 3130 7350 3190
rect 7380 3130 7400 3190
rect 7330 3090 7400 3130
rect 7330 3060 7350 3090
rect 7380 3060 7400 3090
rect 7500 4030 7520 4060
rect 7550 4030 7570 4060
rect 7500 3990 7570 4030
rect 7500 3930 7520 3990
rect 7550 3930 7570 3990
rect 7500 3890 7570 3930
rect 7500 3830 7520 3890
rect 7550 3830 7570 3890
rect 7500 3790 7570 3830
rect 7500 3730 7520 3790
rect 7550 3730 7570 3790
rect 7500 3690 7570 3730
rect 7500 3630 7520 3690
rect 7550 3630 7570 3690
rect 7500 3590 7570 3630
rect 7500 3530 7520 3590
rect 7550 3530 7570 3590
rect 7500 3490 7570 3530
rect 7500 3430 7520 3490
rect 7550 3430 7570 3490
rect 7500 3390 7570 3430
rect 7500 3330 7520 3390
rect 7550 3330 7570 3390
rect 7500 3290 7570 3330
rect 7500 3230 7520 3290
rect 7550 3230 7570 3290
rect 7500 3190 7570 3230
rect 7500 3130 7520 3190
rect 7550 3130 7570 3190
rect 7500 3090 7570 3130
rect 7500 3060 7520 3090
rect 7550 3060 7570 3090
rect 7670 4030 7690 4060
rect 7720 4030 7740 4060
rect 7670 3990 7740 4030
rect 7670 3930 7690 3990
rect 7720 3930 7740 3990
rect 7670 3890 7740 3930
rect 7670 3830 7690 3890
rect 7720 3830 7740 3890
rect 7670 3790 7740 3830
rect 7670 3730 7690 3790
rect 7720 3730 7740 3790
rect 7670 3690 7740 3730
rect 7670 3630 7690 3690
rect 7720 3630 7740 3690
rect 7670 3590 7740 3630
rect 7670 3530 7690 3590
rect 7720 3530 7740 3590
rect 7670 3490 7740 3530
rect 7670 3430 7690 3490
rect 7720 3430 7740 3490
rect 7670 3390 7740 3430
rect 7670 3330 7690 3390
rect 7720 3330 7740 3390
rect 7670 3290 7740 3330
rect 7670 3230 7690 3290
rect 7720 3230 7740 3290
rect 7670 3190 7740 3230
rect 7670 3130 7690 3190
rect 7720 3130 7740 3190
rect 7670 3090 7740 3130
rect 7670 3060 7690 3090
rect 7720 3060 7740 3090
rect 7840 3060 7860 4060
rect 7890 4050 7930 4060
rect 7890 4030 7900 4050
rect 7920 4030 7930 4050
rect 7890 4020 7930 4030
rect 7890 3960 7910 4020
rect 7890 3460 7920 3960
rect 8120 3460 8140 3960
rect 6190 2990 6210 3020
rect 6090 2950 6210 2990
rect 6090 2920 6110 2950
rect 6190 2920 6210 2950
rect 6310 2990 6330 3020
rect 6360 2990 6380 3020
rect 6310 2950 6380 2990
rect 6310 2920 6330 2950
rect 6360 2920 6380 2950
rect 6480 2990 6500 3020
rect 6530 2990 6550 3020
rect 6480 2950 6550 2990
rect 6480 2920 6500 2950
rect 6530 2920 6550 2950
rect 6650 2990 6670 3020
rect 6700 2990 6720 3020
rect 6650 2950 6720 2990
rect 6650 2920 6670 2950
rect 6700 2920 6720 2950
rect 6820 2990 6840 3020
rect 6870 2990 6890 3020
rect 6820 2950 6890 2990
rect 6820 2920 6840 2950
rect 6870 2920 6890 2950
rect 6990 2990 7010 3020
rect 7040 2990 7060 3020
rect 6990 2950 7060 2990
rect 6990 2920 7010 2950
rect 7040 2920 7060 2950
rect 7160 2990 7180 3020
rect 7210 2990 7230 3020
rect 7160 2950 7230 2990
rect 7160 2920 7180 2950
rect 7210 2920 7230 2950
rect 7330 2990 7350 3020
rect 7380 2990 7400 3020
rect 7330 2950 7400 2990
rect 7330 2920 7350 2950
rect 7380 2920 7400 2950
rect 7500 2990 7520 3020
rect 7550 2990 7570 3020
rect 7500 2950 7570 2990
rect 7500 2920 7520 2950
rect 7550 2920 7570 2950
rect 7670 2990 7690 3020
rect 7720 2990 7740 3020
rect 7670 2950 7740 2990
rect 7670 2920 7690 2950
rect 7720 2920 7740 2950
rect 7840 2920 7860 3020
rect 7900 2920 7920 3420
rect 8120 2920 8150 3420
rect 4150 2860 4170 2920
rect 4150 2850 4190 2860
rect 4150 2830 4160 2850
rect 4180 2830 4190 2850
rect 4150 2820 4190 2830
rect 4400 2780 4460 2880
rect 4560 2850 4580 2880
rect 4610 2850 4630 2880
rect 4560 2810 4630 2850
rect 4560 2780 4580 2810
rect 4610 2780 4630 2810
rect 4730 2850 4750 2880
rect 4780 2850 4800 2880
rect 4730 2810 4800 2850
rect 4730 2780 4750 2810
rect 4780 2780 4800 2810
rect 4900 2850 4920 2880
rect 4950 2850 4970 2880
rect 4900 2810 4970 2850
rect 4900 2780 4920 2810
rect 4950 2780 4970 2810
rect 5070 2850 5090 2880
rect 5120 2850 5140 2880
rect 5070 2810 5140 2850
rect 5070 2780 5090 2810
rect 5120 2780 5140 2810
rect 5240 2850 5260 2880
rect 5290 2850 5310 2880
rect 5240 2810 5310 2850
rect 5240 2780 5260 2810
rect 5290 2780 5310 2810
rect 5410 2850 5430 2880
rect 5460 2850 5480 2880
rect 5410 2810 5480 2850
rect 5410 2780 5430 2810
rect 5460 2780 5480 2810
rect 5580 2850 5600 2880
rect 5630 2850 5650 2880
rect 5580 2810 5650 2850
rect 5580 2780 5600 2810
rect 5630 2780 5650 2810
rect 5750 2850 5770 2880
rect 5800 2850 5820 2880
rect 5750 2810 5820 2850
rect 5750 2780 5770 2810
rect 5800 2780 5820 2810
rect 5920 2850 5940 2880
rect 5970 2850 5990 2880
rect 5920 2810 5990 2850
rect 5920 2780 5940 2810
rect 5970 2780 5990 2810
rect 6090 2850 6110 2880
rect 6190 2850 6210 2880
rect 6090 2810 6210 2850
rect 6090 2780 6110 2810
rect 6190 2780 6210 2810
rect 6310 2850 6330 2880
rect 6360 2850 6380 2880
rect 6310 2810 6380 2850
rect 6310 2780 6330 2810
rect 6360 2780 6380 2810
rect 6480 2850 6500 2880
rect 6530 2850 6550 2880
rect 6480 2810 6550 2850
rect 6480 2780 6500 2810
rect 6530 2780 6550 2810
rect 6650 2850 6670 2880
rect 6700 2850 6720 2880
rect 6650 2810 6720 2850
rect 6650 2780 6670 2810
rect 6700 2780 6720 2810
rect 6820 2850 6840 2880
rect 6870 2850 6890 2880
rect 6820 2810 6890 2850
rect 6820 2780 6840 2810
rect 6870 2780 6890 2810
rect 6990 2850 7010 2880
rect 7040 2850 7060 2880
rect 6990 2810 7060 2850
rect 6990 2780 7010 2810
rect 7040 2780 7060 2810
rect 7160 2850 7180 2880
rect 7210 2850 7230 2880
rect 7160 2810 7230 2850
rect 7160 2780 7180 2810
rect 7210 2780 7230 2810
rect 7330 2850 7350 2880
rect 7380 2850 7400 2880
rect 7330 2810 7400 2850
rect 7330 2780 7350 2810
rect 7380 2780 7400 2810
rect 7500 2850 7520 2880
rect 7550 2850 7570 2880
rect 7500 2810 7570 2850
rect 7500 2780 7520 2810
rect 7550 2780 7570 2810
rect 7670 2850 7690 2880
rect 7720 2850 7740 2880
rect 7670 2810 7740 2850
rect 7670 2780 7690 2810
rect 7720 2780 7740 2810
rect 7840 2780 7900 2880
rect 8130 2860 8150 2920
rect 8110 2850 8150 2860
rect 8110 2830 8120 2850
rect 8140 2830 8150 2850
rect 8110 2820 8150 2830
rect 4400 2750 4440 2780
rect 4400 2730 4410 2750
rect 4430 2730 4440 2750
rect 4400 2720 4440 2730
rect 7860 2750 7900 2780
rect 7860 2730 7870 2750
rect 7890 2730 7900 2750
rect 7860 2720 7900 2730
<< polycont >>
rect 4410 7650 4430 7670
rect 7870 7650 7890 7670
rect 4160 7550 4180 7570
rect 8120 7550 8140 7570
rect 4380 6350 4400 6370
rect 7900 6350 7920 6370
rect 4260 6250 4280 6270
rect 4550 6250 4570 6270
rect 4830 6250 4850 6270
rect 5110 6250 5130 6270
rect 5390 6250 5410 6270
rect 5670 6250 5690 6270
rect 6080 6250 6100 6270
rect 6200 6250 6220 6270
rect 6610 6250 6630 6270
rect 6890 6250 6910 6270
rect 7170 6250 7190 6270
rect 7450 6250 7470 6270
rect 7730 6250 7750 6270
rect 8020 6250 8040 6270
rect 4260 4130 4280 4150
rect 4550 4130 4570 4150
rect 4830 4130 4850 4150
rect 5110 4130 5130 4150
rect 5390 4130 5410 4150
rect 5670 4130 5690 4150
rect 6080 4130 6100 4150
rect 6200 4130 6220 4150
rect 6610 4130 6630 4150
rect 6890 4130 6910 4150
rect 7170 4130 7190 4150
rect 7450 4130 7470 4150
rect 7730 4130 7750 4150
rect 8020 4130 8040 4150
rect 4380 4030 4400 4050
rect 7900 4030 7920 4050
rect 4160 2830 4180 2850
rect 8120 2830 8140 2850
rect 4410 2730 4430 2750
rect 7870 2730 7890 2750
<< locali >>
rect 4480 7680 4490 7690
rect 4400 7670 4490 7680
rect 4530 7680 4540 7690
rect 4650 7680 4660 7690
rect 4530 7670 4660 7680
rect 4700 7680 4710 7690
rect 4820 7680 4830 7690
rect 4700 7670 4830 7680
rect 4870 7680 4880 7690
rect 4990 7680 5000 7690
rect 4870 7670 5000 7680
rect 5040 7680 5050 7690
rect 5160 7680 5170 7690
rect 5040 7670 5170 7680
rect 5210 7680 5220 7690
rect 5330 7680 5340 7690
rect 5210 7670 5340 7680
rect 5380 7680 5390 7690
rect 5500 7680 5510 7690
rect 5380 7670 5510 7680
rect 5550 7680 5560 7690
rect 5670 7680 5680 7690
rect 5550 7670 5680 7680
rect 5720 7680 5730 7690
rect 5840 7680 5850 7690
rect 5720 7670 5850 7680
rect 5890 7680 5900 7690
rect 6010 7680 6020 7690
rect 5890 7670 6020 7680
rect 6060 7680 6070 7690
rect 6230 7680 6240 7690
rect 6060 7670 6240 7680
rect 6280 7680 6290 7690
rect 6400 7680 6410 7690
rect 6280 7670 6410 7680
rect 6450 7680 6460 7690
rect 6570 7680 6580 7690
rect 6450 7670 6580 7680
rect 6620 7680 6630 7690
rect 6740 7680 6750 7690
rect 6620 7670 6750 7680
rect 6790 7680 6800 7690
rect 6910 7680 6920 7690
rect 6790 7670 6920 7680
rect 6960 7680 6970 7690
rect 7080 7680 7090 7690
rect 6960 7670 7090 7680
rect 7130 7680 7140 7690
rect 7250 7680 7260 7690
rect 7130 7670 7260 7680
rect 7300 7680 7310 7690
rect 7420 7680 7430 7690
rect 7300 7670 7430 7680
rect 7470 7680 7480 7690
rect 7590 7680 7600 7690
rect 7470 7670 7600 7680
rect 7640 7680 7650 7690
rect 7760 7680 7770 7690
rect 7640 7670 7770 7680
rect 7810 7680 7820 7690
rect 7810 7670 7900 7680
rect 4400 7650 4410 7670
rect 4430 7650 7870 7670
rect 7890 7650 7900 7670
rect 4400 7640 4490 7650
rect 4480 7630 4490 7640
rect 4530 7640 4660 7650
rect 4530 7630 4540 7640
rect 4480 7620 4540 7630
rect 4650 7630 4660 7640
rect 4700 7640 4830 7650
rect 4700 7630 4710 7640
rect 4650 7620 4710 7630
rect 4820 7630 4830 7640
rect 4870 7640 5000 7650
rect 4870 7630 4880 7640
rect 4820 7620 4880 7630
rect 4990 7630 5000 7640
rect 5040 7640 5170 7650
rect 5040 7630 5050 7640
rect 4990 7620 5050 7630
rect 5160 7630 5170 7640
rect 5210 7640 5340 7650
rect 5210 7630 5220 7640
rect 5160 7620 5220 7630
rect 5330 7630 5340 7640
rect 5380 7640 5510 7650
rect 5380 7630 5390 7640
rect 5330 7620 5390 7630
rect 5500 7630 5510 7640
rect 5550 7640 5680 7650
rect 5550 7630 5560 7640
rect 5500 7620 5560 7630
rect 5670 7630 5680 7640
rect 5720 7640 5850 7650
rect 5720 7630 5730 7640
rect 5670 7620 5730 7630
rect 5840 7630 5850 7640
rect 5890 7640 6020 7650
rect 5890 7630 5900 7640
rect 5840 7620 5900 7630
rect 6010 7630 6020 7640
rect 6060 7640 6240 7650
rect 6060 7630 6070 7640
rect 6010 7620 6070 7630
rect 4150 7570 4190 7580
rect 4150 7550 4160 7570
rect 4180 7550 4190 7570
rect 4150 7520 4190 7550
rect 4150 7510 6110 7520
rect 4150 7490 4260 7510
rect 4300 7490 4490 7510
rect 4530 7490 4660 7510
rect 4700 7490 4830 7510
rect 4870 7490 5000 7510
rect 5040 7490 5170 7510
rect 5210 7490 5340 7510
rect 5380 7490 5510 7510
rect 5550 7490 5680 7510
rect 5720 7490 5850 7510
rect 5890 7490 6020 7510
rect 6060 7490 6110 7510
rect 4150 7480 6110 7490
rect 4150 2920 4190 7480
rect 6130 7380 6170 7640
rect 6230 7630 6240 7640
rect 6280 7640 6410 7650
rect 6280 7630 6290 7640
rect 6230 7620 6290 7630
rect 6400 7630 6410 7640
rect 6450 7640 6580 7650
rect 6450 7630 6460 7640
rect 6400 7620 6460 7630
rect 6570 7630 6580 7640
rect 6620 7640 6750 7650
rect 6620 7630 6630 7640
rect 6570 7620 6630 7630
rect 6740 7630 6750 7640
rect 6790 7640 6920 7650
rect 6790 7630 6800 7640
rect 6740 7620 6800 7630
rect 6910 7630 6920 7640
rect 6960 7640 7090 7650
rect 6960 7630 6970 7640
rect 6910 7620 6970 7630
rect 7080 7630 7090 7640
rect 7130 7640 7260 7650
rect 7130 7630 7140 7640
rect 7080 7620 7140 7630
rect 7250 7630 7260 7640
rect 7300 7640 7430 7650
rect 7300 7630 7310 7640
rect 7250 7620 7310 7630
rect 7420 7630 7430 7640
rect 7470 7640 7600 7650
rect 7470 7630 7480 7640
rect 7420 7620 7480 7630
rect 7590 7630 7600 7640
rect 7640 7640 7770 7650
rect 7640 7630 7650 7640
rect 7590 7620 7650 7630
rect 7760 7630 7770 7640
rect 7810 7640 7900 7650
rect 7810 7630 7820 7640
rect 7760 7620 7820 7630
rect 8110 7570 8150 7580
rect 8110 7550 8120 7570
rect 8140 7550 8150 7570
rect 8110 7520 8150 7550
rect 6190 7510 8150 7520
rect 6190 7490 6240 7510
rect 6280 7490 6410 7510
rect 6450 7490 6580 7510
rect 6620 7490 6750 7510
rect 6790 7490 6920 7510
rect 6960 7490 7090 7510
rect 7130 7490 7260 7510
rect 7300 7490 7430 7510
rect 7470 7490 7600 7510
rect 7640 7490 7770 7510
rect 7810 7490 8000 7510
rect 8040 7490 8150 7510
rect 6190 7480 8150 7490
rect 4480 7370 7820 7380
rect 4480 7350 4490 7370
rect 4530 7350 4660 7370
rect 4700 7350 4830 7370
rect 4870 7350 5000 7370
rect 5040 7350 5170 7370
rect 5210 7350 5340 7370
rect 5380 7350 5510 7370
rect 5550 7350 5680 7370
rect 5720 7350 5850 7370
rect 5890 7350 6020 7370
rect 6060 7350 6240 7370
rect 6280 7350 6410 7370
rect 6450 7350 6580 7370
rect 6620 7350 6750 7370
rect 6790 7350 6920 7370
rect 6960 7350 7090 7370
rect 7130 7350 7260 7370
rect 7300 7350 7430 7370
rect 7470 7350 7600 7370
rect 7640 7350 7770 7370
rect 7810 7350 7820 7370
rect 4480 7340 7820 7350
rect 4250 6970 4350 6980
rect 4250 6950 4260 6970
rect 4300 6950 4350 6970
rect 4250 6940 4350 6950
rect 4230 6430 4290 6440
rect 4230 6410 4240 6430
rect 4280 6410 4290 6430
rect 4230 6400 4290 6410
rect 4250 6270 4290 6400
rect 4250 6250 4260 6270
rect 4280 6250 4290 6270
rect 4250 6200 4290 6250
rect 4310 6280 4350 6940
rect 4370 6370 4410 6380
rect 4370 6350 4380 6370
rect 4400 6350 4410 6370
rect 4370 6340 4410 6350
rect 4370 6330 6090 6340
rect 4370 6310 4490 6330
rect 4530 6310 4660 6330
rect 4700 6310 4830 6330
rect 4870 6310 5000 6330
rect 5040 6310 5170 6330
rect 5210 6310 5340 6330
rect 5380 6310 5510 6330
rect 5550 6310 5680 6330
rect 5720 6310 5850 6330
rect 5890 6310 6020 6330
rect 6060 6310 6090 6330
rect 4370 6300 6090 6310
rect 4490 6280 4530 6300
rect 4660 6280 4700 6300
rect 4830 6280 4870 6300
rect 5000 6280 5040 6300
rect 5170 6280 5210 6300
rect 5340 6280 5380 6300
rect 5510 6280 5550 6300
rect 5680 6280 5720 6300
rect 5850 6280 5890 6300
rect 6010 6280 6050 6300
rect 4310 6240 4440 6280
rect 4490 6270 6050 6280
rect 4490 6250 4550 6270
rect 4570 6250 4830 6270
rect 4850 6250 5110 6270
rect 5130 6250 5390 6270
rect 5410 6250 5670 6270
rect 5690 6250 6050 6270
rect 4490 6240 6050 6250
rect 4220 6190 4290 6200
rect 4220 6150 4230 6190
rect 4250 6150 4290 6190
rect 4220 6140 4290 6150
rect 4250 5750 4290 6140
rect 4250 5740 4300 5750
rect 4250 5700 4270 5740
rect 4290 5700 4300 5740
rect 4250 5690 4300 5700
rect 4400 5740 4440 6240
rect 4400 5700 4410 5740
rect 4430 5700 4440 5740
rect 4250 5220 4290 5690
rect 4400 5670 4440 5700
rect 4540 5740 4580 6240
rect 4540 5700 4550 5740
rect 4570 5700 4580 5740
rect 4540 5690 4580 5700
rect 4680 5740 4720 5750
rect 4680 5700 4690 5740
rect 4710 5700 4720 5740
rect 4680 5670 4720 5700
rect 4820 5740 4860 6240
rect 4820 5700 4830 5740
rect 4850 5700 4860 5740
rect 4820 5690 4860 5700
rect 4960 5740 5000 5750
rect 4960 5700 4970 5740
rect 4990 5700 5000 5740
rect 4960 5670 5000 5700
rect 5100 5740 5140 6240
rect 5100 5700 5110 5740
rect 5130 5700 5140 5740
rect 5100 5690 5140 5700
rect 5240 5740 5280 5750
rect 5240 5700 5250 5740
rect 5270 5700 5280 5740
rect 5240 5670 5280 5700
rect 5380 5740 5420 6240
rect 5380 5700 5390 5740
rect 5410 5700 5420 5740
rect 5380 5690 5420 5700
rect 5520 5740 5560 5750
rect 5520 5700 5530 5740
rect 5550 5700 5560 5740
rect 5520 5670 5560 5700
rect 5660 5740 5700 6240
rect 6010 6210 6050 6240
rect 6010 6190 6020 6210
rect 6040 6190 6050 6210
rect 6010 6180 6050 6190
rect 6070 6270 6110 6280
rect 6070 6250 6080 6270
rect 6100 6250 6110 6270
rect 5660 5700 5670 5740
rect 5690 5700 5700 5740
rect 5660 5690 5700 5700
rect 5800 5740 5840 5750
rect 5800 5700 5810 5740
rect 5830 5730 6050 5740
rect 5830 5710 6020 5730
rect 6040 5710 6050 5730
rect 5830 5700 6050 5710
rect 5800 5670 5840 5700
rect 4400 5630 5840 5670
rect 4250 5210 6050 5220
rect 4250 5190 5920 5210
rect 5940 5190 6020 5210
rect 6040 5190 6050 5210
rect 4250 5180 6050 5190
rect 4250 4840 4290 5180
rect 4250 4770 4260 4840
rect 4280 4770 4290 4840
rect 6070 4975 6110 6250
rect 6070 4905 6080 4975
rect 6100 4905 6110 4975
rect 4250 4710 4290 4770
rect 4400 4730 5840 4770
rect 4250 4700 4300 4710
rect 4250 4660 4270 4700
rect 4290 4660 4300 4700
rect 4250 4650 4300 4660
rect 4400 4700 4440 4730
rect 4400 4660 4410 4700
rect 4430 4660 4440 4700
rect 4250 4260 4290 4650
rect 4220 4250 4290 4260
rect 4220 4210 4230 4250
rect 4250 4210 4290 4250
rect 4220 4200 4290 4210
rect 4250 4150 4290 4200
rect 4400 4160 4440 4660
rect 4540 4700 4580 4710
rect 4540 4660 4550 4700
rect 4570 4660 4580 4700
rect 4540 4160 4580 4660
rect 4680 4700 4720 4730
rect 4680 4660 4690 4700
rect 4710 4660 4720 4700
rect 4680 4650 4720 4660
rect 4820 4700 4860 4710
rect 4820 4660 4830 4700
rect 4850 4660 4860 4700
rect 4820 4160 4860 4660
rect 4960 4700 5000 4730
rect 4960 4660 4970 4700
rect 4990 4660 5000 4700
rect 4960 4650 5000 4660
rect 5100 4700 5140 4710
rect 5100 4660 5110 4700
rect 5130 4660 5140 4700
rect 5100 4160 5140 4660
rect 5240 4700 5280 4730
rect 5240 4660 5250 4700
rect 5270 4660 5280 4700
rect 5240 4650 5280 4660
rect 5380 4700 5420 4710
rect 5380 4660 5390 4700
rect 5410 4660 5420 4700
rect 5380 4160 5420 4660
rect 5520 4700 5560 4730
rect 5520 4660 5530 4700
rect 5550 4660 5560 4700
rect 5520 4650 5560 4660
rect 5660 4700 5700 4710
rect 5660 4660 5670 4700
rect 5690 4660 5700 4700
rect 5660 4160 5700 4660
rect 5800 4700 5840 4730
rect 5800 4660 5810 4700
rect 5830 4690 6050 4700
rect 5830 4670 6020 4690
rect 6040 4670 6050 4690
rect 5830 4660 6050 4670
rect 5800 4650 5840 4660
rect 6010 4210 6050 4220
rect 6010 4190 6020 4210
rect 6040 4190 6050 4210
rect 6010 4160 6050 4190
rect 4250 4130 4260 4150
rect 4280 4130 4290 4150
rect 4250 4000 4290 4130
rect 4230 3990 4290 4000
rect 4230 3970 4240 3990
rect 4280 3970 4290 3990
rect 4230 3960 4290 3970
rect 4310 4120 4440 4160
rect 4490 4150 6050 4160
rect 4490 4130 4550 4150
rect 4570 4130 4830 4150
rect 4850 4130 5110 4150
rect 5130 4130 5390 4150
rect 5410 4130 5670 4150
rect 5690 4130 6050 4150
rect 4490 4120 6050 4130
rect 6070 4150 6110 4905
rect 6070 4130 6080 4150
rect 6100 4130 6110 4150
rect 6070 4120 6110 4130
rect 4310 3460 4350 4120
rect 4490 4100 4530 4120
rect 4660 4100 4700 4120
rect 4830 4100 4870 4120
rect 5000 4100 5040 4120
rect 5170 4100 5210 4120
rect 5340 4100 5380 4120
rect 5510 4100 5550 4120
rect 5680 4100 5720 4120
rect 5850 4100 5890 4120
rect 6010 4100 6050 4120
rect 4370 4090 6090 4100
rect 4370 4070 4490 4090
rect 4530 4070 4660 4090
rect 4700 4070 4830 4090
rect 4870 4070 5000 4090
rect 5040 4070 5170 4090
rect 5210 4070 5340 4090
rect 5380 4070 5510 4090
rect 5550 4070 5680 4090
rect 5720 4070 5850 4090
rect 5890 4070 6020 4090
rect 6060 4070 6090 4090
rect 4370 4060 6090 4070
rect 4370 4050 4410 4060
rect 4370 4030 4380 4050
rect 4400 4030 4410 4050
rect 4370 4020 4410 4030
rect 4250 3450 4350 3460
rect 4250 3430 4260 3450
rect 4300 3430 4350 3450
rect 4250 3420 4350 3430
rect 6130 3060 6170 7340
rect 7950 6970 8050 6980
rect 7950 6950 8000 6970
rect 8040 6950 8050 6970
rect 7950 6940 8050 6950
rect 7890 6370 7930 6380
rect 7890 6350 7900 6370
rect 7920 6350 7930 6370
rect 7890 6340 7930 6350
rect 6210 6330 7930 6340
rect 6210 6310 6240 6330
rect 6280 6310 6410 6330
rect 6450 6310 6580 6330
rect 6620 6310 6750 6330
rect 6790 6310 6920 6330
rect 6960 6310 7090 6330
rect 7130 6310 7260 6330
rect 7300 6310 7430 6330
rect 7470 6310 7600 6330
rect 7640 6310 7770 6330
rect 7810 6310 7930 6330
rect 6210 6300 7930 6310
rect 6250 6280 6290 6300
rect 6410 6280 6450 6300
rect 6580 6280 6620 6300
rect 6750 6280 6790 6300
rect 6920 6280 6960 6300
rect 7090 6280 7130 6300
rect 7260 6280 7300 6300
rect 7430 6280 7470 6300
rect 7600 6280 7640 6300
rect 7770 6280 7810 6300
rect 7950 6280 7990 6940
rect 6190 6270 6230 6280
rect 6190 6250 6200 6270
rect 6220 6250 6230 6270
rect 6190 4150 6230 6250
rect 6250 6270 7810 6280
rect 6250 6250 6610 6270
rect 6630 6250 6890 6270
rect 6910 6250 7170 6270
rect 7190 6250 7450 6270
rect 7470 6250 7730 6270
rect 7750 6250 7810 6270
rect 6250 6240 7810 6250
rect 7860 6240 7990 6280
rect 8010 6430 8070 6440
rect 8010 6410 8020 6430
rect 8060 6410 8070 6430
rect 8010 6400 8070 6410
rect 8010 6270 8050 6400
rect 8010 6250 8020 6270
rect 8040 6250 8050 6270
rect 6250 6210 6290 6240
rect 6250 6190 6260 6210
rect 6280 6190 6290 6210
rect 6250 6180 6290 6190
rect 6460 5740 6500 5750
rect 6250 5730 6470 5740
rect 6250 5710 6260 5730
rect 6280 5710 6470 5730
rect 6250 5700 6470 5710
rect 6490 5700 6500 5740
rect 6460 5670 6500 5700
rect 6600 5740 6640 6240
rect 6600 5700 6610 5740
rect 6630 5700 6640 5740
rect 6600 5690 6640 5700
rect 6740 5740 6780 5750
rect 6740 5700 6750 5740
rect 6770 5700 6780 5740
rect 6740 5670 6780 5700
rect 6880 5740 6920 6240
rect 6880 5700 6890 5740
rect 6910 5700 6920 5740
rect 6880 5690 6920 5700
rect 7020 5740 7060 5750
rect 7020 5700 7030 5740
rect 7050 5700 7060 5740
rect 7020 5670 7060 5700
rect 7160 5740 7200 6240
rect 7160 5700 7170 5740
rect 7190 5700 7200 5740
rect 7160 5690 7200 5700
rect 7300 5740 7340 5750
rect 7300 5700 7310 5740
rect 7330 5700 7340 5740
rect 7300 5670 7340 5700
rect 7440 5740 7480 6240
rect 7440 5700 7450 5740
rect 7470 5700 7480 5740
rect 7440 5690 7480 5700
rect 7580 5740 7620 5750
rect 7580 5700 7590 5740
rect 7610 5700 7620 5740
rect 7580 5670 7620 5700
rect 7720 5740 7760 6240
rect 7720 5700 7730 5740
rect 7750 5700 7760 5740
rect 7720 5690 7760 5700
rect 7860 5740 7900 6240
rect 8010 6200 8050 6250
rect 8010 6190 8080 6200
rect 8010 6150 8050 6190
rect 8070 6150 8080 6190
rect 8010 6140 8080 6150
rect 8010 5750 8050 6140
rect 7860 5700 7870 5740
rect 7890 5700 7900 5740
rect 7860 5670 7900 5700
rect 8000 5740 8050 5750
rect 8000 5700 8010 5740
rect 8030 5700 8050 5740
rect 8000 5690 8050 5700
rect 6460 5630 7900 5670
rect 8010 5220 8050 5690
rect 6250 5210 8050 5220
rect 6250 5190 6260 5210
rect 6280 5190 6360 5210
rect 6380 5190 8050 5210
rect 6250 5180 8050 5190
rect 6460 4730 7900 4770
rect 6460 4700 6500 4730
rect 6250 4690 6470 4700
rect 6250 4670 6260 4690
rect 6280 4670 6470 4690
rect 6250 4660 6470 4670
rect 6490 4660 6500 4700
rect 6460 4650 6500 4660
rect 6600 4700 6640 4710
rect 6600 4660 6610 4700
rect 6630 4660 6640 4700
rect 6190 4130 6200 4150
rect 6220 4130 6230 4150
rect 6190 4120 6230 4130
rect 6250 4210 6290 4220
rect 6250 4190 6260 4210
rect 6280 4190 6290 4210
rect 6250 4160 6290 4190
rect 6600 4160 6640 4660
rect 6740 4700 6780 4730
rect 6740 4660 6750 4700
rect 6770 4660 6780 4700
rect 6740 4650 6780 4660
rect 6880 4700 6920 4710
rect 6880 4660 6890 4700
rect 6910 4660 6920 4700
rect 6880 4160 6920 4660
rect 7020 4700 7060 4730
rect 7020 4660 7030 4700
rect 7050 4660 7060 4700
rect 7020 4650 7060 4660
rect 7160 4700 7200 4710
rect 7160 4660 7170 4700
rect 7190 4660 7200 4700
rect 7160 4160 7200 4660
rect 7300 4700 7340 4730
rect 7300 4660 7310 4700
rect 7330 4660 7340 4700
rect 7300 4650 7340 4660
rect 7440 4700 7480 4710
rect 7440 4660 7450 4700
rect 7470 4660 7480 4700
rect 7440 4160 7480 4660
rect 7580 4700 7620 4730
rect 7580 4660 7590 4700
rect 7610 4660 7620 4700
rect 7580 4650 7620 4660
rect 7720 4700 7760 4710
rect 7720 4660 7730 4700
rect 7750 4660 7760 4700
rect 7720 4160 7760 4660
rect 7860 4700 7900 4730
rect 8010 4710 8050 5180
rect 7860 4660 7870 4700
rect 7890 4660 7900 4700
rect 7860 4160 7900 4660
rect 8000 4700 8050 4710
rect 8000 4660 8010 4700
rect 8030 4660 8050 4700
rect 8000 4650 8050 4660
rect 8010 4260 8050 4650
rect 8010 4250 8080 4260
rect 8010 4210 8050 4250
rect 8070 4210 8080 4250
rect 8010 4200 8080 4210
rect 6250 4150 7810 4160
rect 6250 4130 6610 4150
rect 6630 4130 6890 4150
rect 6910 4130 7170 4150
rect 7190 4130 7450 4150
rect 7470 4130 7730 4150
rect 7750 4130 7810 4150
rect 6250 4120 7810 4130
rect 7860 4120 7990 4160
rect 6250 4100 6290 4120
rect 6410 4100 6450 4120
rect 6580 4100 6620 4120
rect 6750 4100 6790 4120
rect 6920 4100 6960 4120
rect 7090 4100 7130 4120
rect 7260 4100 7300 4120
rect 7430 4100 7470 4120
rect 7600 4100 7640 4120
rect 7770 4100 7810 4120
rect 6210 4090 7930 4100
rect 6210 4070 6240 4090
rect 6280 4070 6410 4090
rect 6450 4070 6580 4090
rect 6620 4070 6750 4090
rect 6790 4070 6920 4090
rect 6960 4070 7090 4090
rect 7130 4070 7260 4090
rect 7300 4070 7430 4090
rect 7470 4070 7600 4090
rect 7640 4070 7770 4090
rect 7810 4070 7930 4090
rect 6210 4060 7930 4070
rect 7890 4050 7930 4060
rect 7890 4030 7900 4050
rect 7920 4030 7930 4050
rect 7890 4020 7930 4030
rect 7950 3460 7990 4120
rect 8010 4150 8050 4200
rect 8010 4130 8020 4150
rect 8040 4130 8050 4150
rect 8010 4000 8050 4130
rect 8010 3990 8070 4000
rect 8010 3970 8020 3990
rect 8060 3970 8070 3990
rect 8010 3960 8070 3970
rect 7950 3450 8050 3460
rect 7950 3430 8000 3450
rect 8040 3430 8050 3450
rect 7950 3420 8050 3430
rect 4480 3050 7820 3060
rect 4480 3030 4490 3050
rect 4530 3030 4660 3050
rect 4700 3030 4830 3050
rect 4870 3030 5000 3050
rect 5040 3030 5170 3050
rect 5210 3030 5340 3050
rect 5380 3030 5510 3050
rect 5550 3030 5680 3050
rect 5720 3030 5850 3050
rect 5890 3030 6020 3050
rect 6060 3030 6240 3050
rect 6280 3030 6410 3050
rect 6450 3030 6580 3050
rect 6620 3030 6750 3050
rect 6790 3030 6920 3050
rect 6960 3030 7090 3050
rect 7130 3030 7260 3050
rect 7300 3030 7430 3050
rect 7470 3030 7600 3050
rect 7640 3030 7770 3050
rect 7810 3030 7820 3050
rect 4480 3020 7820 3030
rect 4150 2910 6110 2920
rect 4150 2890 4260 2910
rect 4300 2890 4490 2910
rect 4530 2890 4660 2910
rect 4700 2890 4830 2910
rect 4870 2890 5000 2910
rect 5040 2890 5170 2910
rect 5210 2890 5340 2910
rect 5380 2890 5510 2910
rect 5550 2890 5680 2910
rect 5720 2890 5850 2910
rect 5890 2890 6020 2910
rect 6060 2890 6110 2910
rect 4150 2880 6110 2890
rect 4150 2855 4190 2880
rect 4120 2850 4190 2855
rect 4120 2830 4160 2850
rect 4180 2830 4190 2850
rect 4120 2820 4190 2830
rect 4480 2770 4540 2780
rect 4480 2760 4490 2770
rect 4150 2750 4490 2760
rect 4530 2760 4540 2770
rect 4650 2770 4710 2780
rect 4650 2760 4660 2770
rect 4530 2750 4660 2760
rect 4700 2760 4710 2770
rect 4820 2770 4880 2780
rect 4820 2760 4830 2770
rect 4700 2750 4830 2760
rect 4870 2760 4880 2770
rect 4990 2770 5050 2780
rect 4990 2760 5000 2770
rect 4870 2750 5000 2760
rect 5040 2760 5050 2770
rect 5160 2770 5220 2780
rect 5160 2760 5170 2770
rect 5040 2750 5170 2760
rect 5210 2760 5220 2770
rect 5330 2770 5390 2780
rect 5330 2760 5340 2770
rect 5210 2750 5340 2760
rect 5380 2760 5390 2770
rect 5500 2770 5560 2780
rect 5500 2760 5510 2770
rect 5380 2750 5510 2760
rect 5550 2760 5560 2770
rect 5670 2770 5730 2780
rect 5670 2760 5680 2770
rect 5550 2750 5680 2760
rect 5720 2760 5730 2770
rect 5840 2770 5900 2780
rect 5840 2760 5850 2770
rect 5720 2750 5850 2760
rect 5890 2760 5900 2770
rect 6010 2770 6070 2780
rect 6010 2760 6020 2770
rect 5890 2750 6020 2760
rect 6060 2760 6070 2770
rect 6130 2760 6170 3020
rect 8110 2920 8150 7480
rect 6190 2910 8150 2920
rect 6190 2890 6240 2910
rect 6280 2890 6410 2910
rect 6450 2890 6580 2910
rect 6620 2890 6750 2910
rect 6790 2890 6920 2910
rect 6960 2890 7090 2910
rect 7130 2890 7260 2910
rect 7300 2890 7430 2910
rect 7470 2890 7600 2910
rect 7640 2890 7770 2910
rect 7810 2890 8000 2910
rect 8040 2890 8150 2910
rect 6190 2880 8150 2890
rect 8110 2850 8150 2880
rect 8110 2830 8120 2850
rect 8140 2830 8150 2850
rect 8110 2820 8150 2830
rect 6230 2770 6290 2780
rect 6230 2760 6240 2770
rect 6060 2750 6240 2760
rect 6280 2760 6290 2770
rect 6400 2770 6460 2780
rect 6400 2760 6410 2770
rect 6280 2750 6410 2760
rect 6450 2760 6460 2770
rect 6570 2770 6630 2780
rect 6570 2760 6580 2770
rect 6450 2750 6580 2760
rect 6620 2760 6630 2770
rect 6740 2770 6800 2780
rect 6740 2760 6750 2770
rect 6620 2750 6750 2760
rect 6790 2760 6800 2770
rect 6910 2770 6970 2780
rect 6910 2760 6920 2770
rect 6790 2750 6920 2760
rect 6960 2760 6970 2770
rect 7080 2770 7140 2780
rect 7080 2760 7090 2770
rect 6960 2750 7090 2760
rect 7130 2760 7140 2770
rect 7250 2770 7310 2780
rect 7250 2760 7260 2770
rect 7130 2750 7260 2760
rect 7300 2760 7310 2770
rect 7420 2770 7480 2780
rect 7420 2760 7430 2770
rect 7300 2750 7430 2760
rect 7470 2760 7480 2770
rect 7590 2770 7650 2780
rect 7590 2760 7600 2770
rect 7470 2750 7600 2760
rect 7640 2760 7650 2770
rect 7760 2770 7820 2780
rect 7760 2760 7770 2770
rect 7640 2750 7770 2760
rect 7810 2760 7820 2770
rect 7810 2750 8150 2760
rect 4150 2730 4410 2750
rect 4430 2730 7870 2750
rect 7890 2730 8150 2750
rect 4150 2720 4490 2730
rect 4480 2710 4490 2720
rect 4530 2720 4660 2730
rect 4530 2710 4540 2720
rect 4650 2710 4660 2720
rect 4700 2720 4830 2730
rect 4700 2710 4710 2720
rect 4820 2710 4830 2720
rect 4870 2720 5000 2730
rect 4870 2710 4880 2720
rect 4990 2710 5000 2720
rect 5040 2720 5170 2730
rect 5040 2710 5050 2720
rect 5160 2710 5170 2720
rect 5210 2720 5340 2730
rect 5210 2710 5220 2720
rect 5330 2710 5340 2720
rect 5380 2720 5510 2730
rect 5380 2710 5390 2720
rect 5500 2710 5510 2720
rect 5550 2720 5680 2730
rect 5550 2710 5560 2720
rect 5670 2710 5680 2720
rect 5720 2720 5850 2730
rect 5720 2710 5730 2720
rect 5840 2710 5850 2720
rect 5890 2720 6020 2730
rect 5890 2710 5900 2720
rect 6010 2710 6020 2720
rect 6060 2720 6240 2730
rect 6060 2710 6070 2720
rect 6230 2710 6240 2720
rect 6280 2720 6410 2730
rect 6280 2710 6290 2720
rect 6400 2710 6410 2720
rect 6450 2720 6580 2730
rect 6450 2710 6460 2720
rect 6570 2710 6580 2720
rect 6620 2720 6750 2730
rect 6620 2710 6630 2720
rect 6740 2710 6750 2720
rect 6790 2720 6920 2730
rect 6790 2710 6800 2720
rect 6910 2710 6920 2720
rect 6960 2720 7090 2730
rect 6960 2710 6970 2720
rect 7080 2710 7090 2720
rect 7130 2720 7260 2730
rect 7130 2710 7140 2720
rect 7250 2710 7260 2720
rect 7300 2720 7430 2730
rect 7300 2710 7310 2720
rect 7420 2710 7430 2720
rect 7470 2720 7600 2730
rect 7470 2710 7480 2720
rect 7590 2710 7600 2720
rect 7640 2720 7770 2730
rect 7640 2710 7650 2720
rect 7760 2710 7770 2720
rect 7810 2720 8150 2730
rect 7810 2710 7820 2720
<< viali >>
rect 4260 4770 4280 4840
rect 6080 4905 6100 4975
<< metal1 >>
rect 4115 4975 6110 4985
rect 4115 4905 6080 4975
rect 6100 4905 6110 4975
rect 4115 4895 6110 4905
rect 4115 4840 4290 4850
rect 4115 4770 4260 4840
rect 4280 4770 4290 4840
rect 4115 4760 4290 4770
<< labels >>
rlabel locali 4150 2740 4150 2740 7 VN
port 1 w
rlabel metal1 4115 4935 4115 4935 7 Vbn
port 2 w
rlabel locali 4120 2835 4120 2835 7 Vc
port 3 w
rlabel metal1 4115 4805 4115 4805 7 VP
port 4 w
<< end >>
