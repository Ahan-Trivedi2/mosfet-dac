magic
tech sky130A
timestamp 1762137910
<< nwell >>
rect -20 4400 3400 5830
rect -20 810 3400 2240
<< nmos >>
rect -280 5100 -80 5600
rect -280 4560 -80 5060
rect 3460 5100 3660 5600
rect 3460 4560 3660 5060
rect -160 3340 -60 4340
rect -20 3340 80 4340
rect 120 3340 220 4340
rect 260 3340 360 4340
rect 400 3340 500 4340
rect 540 3340 640 4340
rect 680 3340 780 4340
rect 820 3340 920 4340
rect 960 3340 1060 4340
rect 1100 3340 1200 4340
rect 1240 3340 1340 4340
rect -160 2300 -60 3300
rect -20 2300 80 3300
rect 120 2300 220 3300
rect 260 2300 360 3300
rect 400 2300 500 3300
rect 540 2300 640 3300
rect 680 2300 780 3300
rect 820 2300 920 3300
rect 960 2300 1060 3300
rect 1100 2300 1200 3300
rect 1240 2300 1340 3300
rect 2040 3340 2140 4340
rect 2180 3340 2280 4340
rect 2320 3340 2420 4340
rect 2460 3340 2560 4340
rect 2600 3340 2700 4340
rect 2740 3340 2840 4340
rect 2880 3340 2980 4340
rect 3020 3340 3120 4340
rect 3160 3340 3260 4340
rect 3300 3340 3400 4340
rect 3440 3340 3540 4340
rect 2040 2300 2140 3300
rect 2180 2300 2280 3300
rect 2320 2300 2420 3300
rect 2460 2300 2560 3300
rect 2600 2300 2700 3300
rect 2740 2300 2840 3300
rect 2880 2300 2980 3300
rect 3020 2300 3120 3300
rect 3160 2300 3260 3300
rect 3300 2300 3400 3300
rect 3440 2300 3540 3300
rect -280 1580 -80 2080
rect -280 1040 -80 1540
rect 3460 1580 3660 2080
rect 3460 1040 3660 1540
<< pmos >>
rect 0 5640 100 5740
rect 170 5640 270 5740
rect 340 5640 440 5740
rect 510 5640 610 5740
rect 680 5640 780 5740
rect 850 5640 950 5740
rect 1020 5640 1120 5740
rect 1190 5640 1290 5740
rect 1360 5640 1460 5740
rect 1530 5640 1630 5740
rect 1750 5640 1850 5740
rect 1920 5640 2020 5740
rect 2090 5640 2190 5740
rect 2260 5640 2360 5740
rect 2430 5640 2530 5740
rect 2600 5640 2700 5740
rect 2770 5640 2870 5740
rect 2940 5640 3040 5740
rect 3110 5640 3210 5740
rect 3280 5640 3380 5740
rect 0 5500 100 5600
rect 170 5500 270 5600
rect 340 5500 440 5600
rect 510 5500 610 5600
rect 680 5500 780 5600
rect 850 5500 950 5600
rect 1020 5500 1120 5600
rect 1190 5500 1290 5600
rect 1360 5500 1460 5600
rect 1530 5500 1630 5600
rect 0 4460 100 5460
rect 170 4460 270 5460
rect 340 4460 440 5460
rect 510 4460 610 5460
rect 680 4460 780 5460
rect 850 4460 950 5460
rect 1020 4460 1120 5460
rect 1190 4460 1290 5460
rect 1360 4460 1460 5460
rect 1530 4460 1630 5460
rect 1750 5500 1850 5600
rect 1920 5500 2020 5600
rect 2090 5500 2190 5600
rect 2260 5500 2360 5600
rect 2430 5500 2530 5600
rect 2600 5500 2700 5600
rect 2770 5500 2870 5600
rect 2940 5500 3040 5600
rect 3110 5500 3210 5600
rect 3280 5500 3380 5600
rect 1750 4460 1850 5460
rect 1920 4460 2020 5460
rect 2090 4460 2190 5460
rect 2260 4460 2360 5460
rect 2430 4460 2530 5460
rect 2600 4460 2700 5460
rect 2770 4460 2870 5460
rect 2940 4460 3040 5460
rect 3110 4460 3210 5460
rect 3280 4460 3380 5460
rect 0 1180 100 2180
rect 170 1180 270 2180
rect 340 1180 440 2180
rect 510 1180 610 2180
rect 680 1180 780 2180
rect 850 1180 950 2180
rect 1020 1180 1120 2180
rect 1190 1180 1290 2180
rect 1360 1180 1460 2180
rect 1530 1180 1630 2180
rect 0 1040 100 1140
rect 170 1040 270 1140
rect 340 1040 440 1140
rect 510 1040 610 1140
rect 680 1040 780 1140
rect 850 1040 950 1140
rect 1020 1040 1120 1140
rect 1190 1040 1290 1140
rect 1360 1040 1460 1140
rect 1530 1040 1630 1140
rect 1750 1180 1850 2180
rect 1920 1180 2020 2180
rect 2090 1180 2190 2180
rect 2260 1180 2360 2180
rect 2430 1180 2530 2180
rect 2600 1180 2700 2180
rect 2770 1180 2870 2180
rect 2940 1180 3040 2180
rect 3110 1180 3210 2180
rect 3280 1180 3380 2180
rect 1750 1040 1850 1140
rect 1920 1040 2020 1140
rect 2090 1040 2190 1140
rect 2260 1040 2360 1140
rect 2430 1040 2530 1140
rect 2600 1040 2700 1140
rect 2770 1040 2870 1140
rect 2940 1040 3040 1140
rect 3110 1040 3210 1140
rect 3280 1040 3380 1140
rect 0 900 100 1000
rect 170 900 270 1000
rect 340 900 440 1000
rect 510 900 610 1000
rect 680 900 780 1000
rect 850 900 950 1000
rect 1020 900 1120 1000
rect 1190 900 1290 1000
rect 1360 900 1460 1000
rect 1530 900 1630 1000
rect 1750 900 1850 1000
rect 1920 900 2020 1000
rect 2090 900 2190 1000
rect 2260 900 2360 1000
rect 2430 900 2530 1000
rect 2600 900 2700 1000
rect 2770 900 2870 1000
rect 2940 900 3040 1000
rect 3110 900 3210 1000
rect 3280 900 3380 1000
<< ndiff >>
rect -280 5630 -80 5640
rect -280 5610 -200 5630
rect -160 5610 -80 5630
rect -280 5600 -80 5610
rect 3460 5630 3660 5640
rect 3460 5610 3540 5630
rect 3580 5610 3660 5630
rect 3460 5600 3660 5610
rect -280 5090 -80 5100
rect -280 5070 -200 5090
rect -160 5070 -80 5090
rect -280 5060 -80 5070
rect -280 4550 -80 4560
rect -280 4530 -220 4550
rect -180 4530 -80 4550
rect -280 4520 -80 4530
rect 3460 5090 3660 5100
rect 3460 5070 3540 5090
rect 3580 5070 3660 5090
rect 3460 5060 3660 5070
rect 3460 4550 3660 4560
rect 3460 4530 3560 4550
rect 3600 4530 3660 4550
rect 3460 4520 3660 4530
rect -240 4320 -160 4340
rect -200 4260 -160 4320
rect -240 3860 -160 4260
rect -240 3820 -190 3860
rect -170 3820 -160 3860
rect -240 3340 -160 3820
rect -60 3860 -20 4340
rect -60 3820 -50 3860
rect -30 3820 -20 3860
rect -60 3340 -20 3820
rect 80 3860 120 4340
rect 80 3820 90 3860
rect 110 3820 120 3860
rect 80 3340 120 3820
rect 220 3860 260 4340
rect 220 3820 230 3860
rect 250 3820 260 3860
rect 220 3340 260 3820
rect 360 3860 400 4340
rect 360 3820 370 3860
rect 390 3820 400 3860
rect 360 3340 400 3820
rect 500 3860 540 4340
rect 500 3820 510 3860
rect 530 3820 540 3860
rect 500 3340 540 3820
rect 640 3860 680 4340
rect 640 3820 650 3860
rect 670 3820 680 3860
rect 640 3340 680 3820
rect 780 3860 820 4340
rect 780 3820 790 3860
rect 810 3820 820 3860
rect 780 3340 820 3820
rect 920 3860 960 4340
rect 920 3820 930 3860
rect 950 3820 960 3860
rect 920 3340 960 3820
rect 1060 3860 1100 4340
rect 1060 3820 1070 3860
rect 1090 3820 1100 3860
rect 1060 3340 1100 3820
rect 1200 3860 1240 4340
rect 1200 3820 1210 3860
rect 1230 3820 1240 3860
rect 1200 3340 1240 3820
rect 1340 3860 1380 4340
rect 1550 4330 1830 4340
rect 1550 4310 1560 4330
rect 1580 4310 1800 4330
rect 1820 4310 1830 4330
rect 1550 4300 1830 4310
rect 2000 3860 2040 4340
rect 1340 3820 1350 3860
rect 1370 3820 1380 3860
rect 1550 3850 1830 3860
rect 1550 3830 1560 3850
rect 1580 3830 1800 3850
rect 1820 3830 1830 3850
rect 1550 3820 1830 3830
rect 2000 3820 2010 3860
rect 2030 3820 2040 3860
rect 1340 3340 1380 3820
rect -240 3300 -170 3340
rect -50 3300 -30 3340
rect 90 3300 110 3340
rect 230 3300 250 3340
rect 370 3300 390 3340
rect 510 3300 530 3340
rect 650 3300 670 3340
rect 790 3300 810 3340
rect 930 3300 950 3340
rect 1070 3300 1090 3340
rect 1210 3300 1230 3340
rect 1350 3300 1370 3340
rect -240 2820 -160 3300
rect -240 2780 -190 2820
rect -170 2780 -160 2820
rect -240 2380 -160 2780
rect -200 2320 -160 2380
rect -240 2300 -160 2320
rect -60 2820 -20 3300
rect -60 2780 -50 2820
rect -30 2780 -20 2820
rect -60 2300 -20 2780
rect 80 2820 120 3300
rect 80 2780 90 2820
rect 110 2780 120 2820
rect 80 2300 120 2780
rect 220 2820 260 3300
rect 220 2780 230 2820
rect 250 2780 260 2820
rect 220 2300 260 2780
rect 360 2820 400 3300
rect 360 2780 370 2820
rect 390 2780 400 2820
rect 360 2300 400 2780
rect 500 2820 540 3300
rect 500 2780 510 2820
rect 530 2780 540 2820
rect 500 2300 540 2780
rect 640 2820 680 3300
rect 640 2780 650 2820
rect 670 2780 680 2820
rect 640 2300 680 2780
rect 780 2820 820 3300
rect 780 2780 790 2820
rect 810 2780 820 2820
rect 780 2300 820 2780
rect 920 2820 960 3300
rect 920 2780 930 2820
rect 950 2780 960 2820
rect 920 2300 960 2780
rect 1060 2820 1100 3300
rect 1060 2780 1070 2820
rect 1090 2780 1100 2820
rect 1060 2300 1100 2780
rect 1200 2820 1240 3300
rect 1200 2780 1210 2820
rect 1230 2780 1240 2820
rect 1200 2300 1240 2780
rect 1340 2820 1380 3300
rect 1550 3330 1830 3340
rect 1550 3310 1560 3330
rect 1580 3310 1800 3330
rect 1820 3310 1830 3330
rect 1550 3300 1830 3310
rect 2000 3340 2040 3820
rect 2140 3860 2180 4340
rect 2140 3820 2150 3860
rect 2170 3820 2180 3860
rect 2140 3340 2180 3820
rect 2280 3860 2320 4340
rect 2280 3820 2290 3860
rect 2310 3820 2320 3860
rect 2280 3340 2320 3820
rect 2420 3860 2460 4340
rect 2420 3820 2430 3860
rect 2450 3820 2460 3860
rect 2420 3340 2460 3820
rect 2560 3860 2600 4340
rect 2560 3820 2570 3860
rect 2590 3820 2600 3860
rect 2560 3340 2600 3820
rect 2700 3860 2740 4340
rect 2700 3820 2710 3860
rect 2730 3820 2740 3860
rect 2700 3340 2740 3820
rect 2840 3860 2880 4340
rect 2840 3820 2850 3860
rect 2870 3820 2880 3860
rect 2840 3340 2880 3820
rect 2980 3860 3020 4340
rect 2980 3820 2990 3860
rect 3010 3820 3020 3860
rect 2980 3340 3020 3820
rect 3120 3860 3160 4340
rect 3120 3820 3130 3860
rect 3150 3820 3160 3860
rect 3120 3340 3160 3820
rect 3260 3860 3300 4340
rect 3260 3820 3270 3860
rect 3290 3820 3300 3860
rect 3260 3340 3300 3820
rect 3400 3860 3440 4340
rect 3400 3820 3410 3860
rect 3430 3820 3440 3860
rect 3400 3340 3440 3820
rect 3540 4320 3620 4340
rect 3540 4260 3580 4320
rect 3540 3860 3620 4260
rect 3540 3820 3550 3860
rect 3570 3820 3620 3860
rect 3540 3340 3620 3820
rect 2010 3300 2030 3340
rect 2150 3300 2170 3340
rect 2290 3300 2310 3340
rect 2430 3300 2450 3340
rect 2570 3300 2590 3340
rect 2710 3300 2730 3340
rect 2850 3300 2870 3340
rect 2990 3300 3010 3340
rect 3130 3300 3150 3340
rect 3270 3300 3290 3340
rect 3410 3300 3430 3340
rect 3550 3300 3620 3340
rect 2000 2820 2040 3300
rect 1340 2780 1350 2820
rect 1370 2780 1380 2820
rect 1550 2810 1830 2820
rect 1550 2790 1560 2810
rect 1580 2790 1800 2810
rect 1820 2790 1830 2810
rect 1550 2780 1830 2790
rect 2000 2780 2010 2820
rect 2030 2780 2040 2820
rect 1340 2300 1380 2780
rect 1550 2330 1830 2340
rect 1550 2310 1560 2330
rect 1580 2310 1800 2330
rect 1820 2310 1830 2330
rect 1550 2300 1830 2310
rect 2000 2300 2040 2780
rect 2140 2820 2180 3300
rect 2140 2780 2150 2820
rect 2170 2780 2180 2820
rect 2140 2300 2180 2780
rect 2280 2820 2320 3300
rect 2280 2780 2290 2820
rect 2310 2780 2320 2820
rect 2280 2300 2320 2780
rect 2420 2820 2460 3300
rect 2420 2780 2430 2820
rect 2450 2780 2460 2820
rect 2420 2300 2460 2780
rect 2560 2820 2600 3300
rect 2560 2780 2570 2820
rect 2590 2780 2600 2820
rect 2560 2300 2600 2780
rect 2700 2820 2740 3300
rect 2700 2780 2710 2820
rect 2730 2780 2740 2820
rect 2700 2300 2740 2780
rect 2840 2820 2880 3300
rect 2840 2780 2850 2820
rect 2870 2780 2880 2820
rect 2840 2300 2880 2780
rect 2980 2820 3020 3300
rect 2980 2780 2990 2820
rect 3010 2780 3020 2820
rect 2980 2300 3020 2780
rect 3120 2820 3160 3300
rect 3120 2780 3130 2820
rect 3150 2780 3160 2820
rect 3120 2300 3160 2780
rect 3260 2820 3300 3300
rect 3260 2780 3270 2820
rect 3290 2780 3300 2820
rect 3260 2300 3300 2780
rect 3400 2820 3440 3300
rect 3400 2780 3410 2820
rect 3430 2780 3440 2820
rect 3400 2300 3440 2780
rect 3540 2820 3620 3300
rect 3540 2780 3550 2820
rect 3570 2780 3620 2820
rect 3540 2380 3620 2780
rect 3540 2320 3580 2380
rect 3540 2300 3620 2320
rect -280 2110 -80 2120
rect -280 2090 -220 2110
rect -180 2090 -80 2110
rect -280 2080 -80 2090
rect -280 1570 -80 1580
rect -280 1550 -200 1570
rect -160 1550 -80 1570
rect -280 1540 -80 1550
rect 3460 2110 3660 2120
rect 3460 2090 3560 2110
rect 3600 2090 3660 2110
rect 3460 2080 3660 2090
rect 3460 1570 3660 1580
rect 3460 1550 3540 1570
rect 3580 1550 3660 1570
rect 3460 1540 3660 1550
rect -280 1030 -80 1040
rect -280 1010 -200 1030
rect -160 1010 -80 1030
rect -280 1000 -80 1010
rect 3460 1030 3660 1040
rect 3460 1010 3540 1030
rect 3580 1010 3660 1030
rect 3460 1000 3660 1010
<< pdiff >>
rect 0 5770 100 5780
rect 0 5750 30 5770
rect 70 5750 100 5770
rect 0 5740 100 5750
rect 170 5770 270 5780
rect 170 5750 200 5770
rect 240 5750 270 5770
rect 170 5740 270 5750
rect 340 5770 440 5780
rect 340 5750 370 5770
rect 410 5750 440 5770
rect 340 5740 440 5750
rect 510 5770 610 5780
rect 510 5750 540 5770
rect 580 5750 610 5770
rect 510 5740 610 5750
rect 680 5770 780 5780
rect 680 5750 710 5770
rect 750 5750 780 5770
rect 680 5740 780 5750
rect 850 5770 950 5780
rect 850 5750 880 5770
rect 920 5750 950 5770
rect 850 5740 950 5750
rect 1020 5770 1120 5780
rect 1020 5750 1050 5770
rect 1090 5750 1120 5770
rect 1020 5740 1120 5750
rect 1190 5770 1290 5780
rect 1190 5750 1220 5770
rect 1260 5750 1290 5770
rect 1190 5740 1290 5750
rect 1360 5770 1460 5780
rect 1360 5750 1390 5770
rect 1430 5750 1460 5770
rect 1360 5740 1460 5750
rect 1530 5770 1630 5780
rect 1530 5750 1560 5770
rect 1600 5750 1630 5770
rect 1530 5740 1630 5750
rect 1750 5770 1850 5780
rect 1750 5750 1780 5770
rect 1820 5750 1850 5770
rect 1750 5740 1850 5750
rect 1920 5770 2020 5780
rect 1920 5750 1950 5770
rect 1990 5750 2020 5770
rect 1920 5740 2020 5750
rect 2090 5770 2190 5780
rect 2090 5750 2120 5770
rect 2160 5750 2190 5770
rect 2090 5740 2190 5750
rect 2260 5770 2360 5780
rect 2260 5750 2290 5770
rect 2330 5750 2360 5770
rect 2260 5740 2360 5750
rect 2430 5770 2530 5780
rect 2430 5750 2460 5770
rect 2500 5750 2530 5770
rect 2430 5740 2530 5750
rect 2600 5770 2700 5780
rect 2600 5750 2630 5770
rect 2670 5750 2700 5770
rect 2600 5740 2700 5750
rect 2770 5770 2870 5780
rect 2770 5750 2800 5770
rect 2840 5750 2870 5770
rect 2770 5740 2870 5750
rect 2940 5770 3040 5780
rect 2940 5750 2970 5770
rect 3010 5750 3040 5770
rect 2940 5740 3040 5750
rect 3110 5770 3210 5780
rect 3110 5750 3140 5770
rect 3180 5750 3210 5770
rect 3110 5740 3210 5750
rect 3280 5770 3380 5780
rect 3280 5750 3310 5770
rect 3350 5750 3380 5770
rect 3280 5740 3380 5750
rect 0 5630 100 5640
rect 170 5630 270 5640
rect 340 5630 440 5640
rect 510 5630 610 5640
rect 680 5630 780 5640
rect 850 5630 950 5640
rect 1020 5630 1120 5640
rect 1190 5630 1290 5640
rect 1360 5630 1460 5640
rect 1530 5630 1630 5640
rect 1750 5630 1850 5640
rect 1920 5630 2020 5640
rect 2090 5630 2190 5640
rect 2260 5630 2360 5640
rect 2430 5630 2530 5640
rect 2600 5630 2700 5640
rect 2770 5630 2870 5640
rect 2940 5630 3040 5640
rect 3110 5630 3210 5640
rect 3280 5630 3380 5640
rect 0 5610 30 5630
rect 70 5610 200 5630
rect 240 5610 370 5630
rect 410 5610 540 5630
rect 580 5610 710 5630
rect 750 5610 880 5630
rect 920 5610 1050 5630
rect 1090 5610 1220 5630
rect 1260 5610 1390 5630
rect 1430 5610 1560 5630
rect 1600 5610 1780 5630
rect 1820 5610 1950 5630
rect 1990 5610 2120 5630
rect 2160 5610 2290 5630
rect 2330 5610 2460 5630
rect 2500 5610 2630 5630
rect 2670 5610 2800 5630
rect 2840 5610 2970 5630
rect 3010 5610 3140 5630
rect 3180 5610 3310 5630
rect 3350 5610 3380 5630
rect 0 5600 100 5610
rect 170 5600 270 5610
rect 340 5600 440 5610
rect 510 5600 610 5610
rect 680 5600 780 5610
rect 850 5600 950 5610
rect 1020 5600 1120 5610
rect 1190 5600 1290 5610
rect 1360 5600 1460 5610
rect 1530 5600 1630 5610
rect 1750 5600 1850 5610
rect 1920 5600 2020 5610
rect 2090 5600 2190 5610
rect 2260 5600 2360 5610
rect 2430 5600 2530 5610
rect 2600 5600 2700 5610
rect 2770 5600 2870 5610
rect 2940 5600 3040 5610
rect 3110 5600 3210 5610
rect 3280 5600 3380 5610
rect 0 5490 100 5500
rect 0 5470 30 5490
rect 70 5470 100 5490
rect 0 5460 100 5470
rect 170 5490 270 5500
rect 170 5470 200 5490
rect 240 5470 270 5490
rect 170 5460 270 5470
rect 340 5490 440 5500
rect 340 5470 370 5490
rect 410 5470 440 5490
rect 340 5460 440 5470
rect 510 5490 610 5500
rect 510 5470 540 5490
rect 580 5470 610 5490
rect 510 5460 610 5470
rect 680 5490 780 5500
rect 680 5470 710 5490
rect 750 5470 780 5490
rect 680 5460 780 5470
rect 850 5490 950 5500
rect 850 5470 880 5490
rect 920 5470 950 5490
rect 850 5460 950 5470
rect 1020 5490 1120 5500
rect 1020 5470 1050 5490
rect 1090 5470 1120 5490
rect 1020 5460 1120 5470
rect 1190 5490 1290 5500
rect 1190 5470 1220 5490
rect 1260 5470 1290 5490
rect 1190 5460 1290 5470
rect 1360 5490 1460 5500
rect 1360 5470 1390 5490
rect 1430 5470 1460 5490
rect 1360 5460 1460 5470
rect 1530 5490 1630 5500
rect 1530 5470 1560 5490
rect 1600 5470 1630 5490
rect 1530 5460 1630 5470
rect 1750 5490 1850 5500
rect 1750 5470 1780 5490
rect 1820 5470 1850 5490
rect 1750 5460 1850 5470
rect 1920 5490 2020 5500
rect 1920 5470 1950 5490
rect 1990 5470 2020 5490
rect 1920 5460 2020 5470
rect 2090 5490 2190 5500
rect 2090 5470 2120 5490
rect 2160 5470 2190 5490
rect 2090 5460 2190 5470
rect 2260 5490 2360 5500
rect 2260 5470 2290 5490
rect 2330 5470 2360 5490
rect 2260 5460 2360 5470
rect 2430 5490 2530 5500
rect 2430 5470 2460 5490
rect 2500 5470 2530 5490
rect 2430 5460 2530 5470
rect 2600 5490 2700 5500
rect 2600 5470 2630 5490
rect 2670 5470 2700 5490
rect 2600 5460 2700 5470
rect 2770 5490 2870 5500
rect 2770 5470 2800 5490
rect 2840 5470 2870 5490
rect 2770 5460 2870 5470
rect 2940 5490 3040 5500
rect 2940 5470 2970 5490
rect 3010 5470 3040 5490
rect 2940 5460 3040 5470
rect 3110 5490 3210 5500
rect 3110 5470 3140 5490
rect 3180 5470 3210 5490
rect 3110 5460 3210 5470
rect 3280 5490 3380 5500
rect 3280 5470 3310 5490
rect 3350 5470 3380 5490
rect 3280 5460 3380 5470
rect 0 4450 100 4460
rect 0 4430 30 4450
rect 70 4430 100 4450
rect 0 4420 100 4430
rect 170 4450 270 4460
rect 170 4430 200 4450
rect 240 4430 270 4450
rect 170 4420 270 4430
rect 340 4450 440 4460
rect 340 4430 370 4450
rect 410 4430 440 4450
rect 340 4420 440 4430
rect 510 4450 610 4460
rect 510 4430 540 4450
rect 580 4430 610 4450
rect 510 4420 610 4430
rect 680 4450 780 4460
rect 680 4430 710 4450
rect 750 4430 780 4450
rect 680 4420 780 4430
rect 850 4450 950 4460
rect 850 4430 880 4450
rect 920 4430 950 4450
rect 850 4420 950 4430
rect 1020 4450 1120 4460
rect 1020 4430 1050 4450
rect 1090 4430 1120 4450
rect 1020 4420 1120 4430
rect 1190 4450 1290 4460
rect 1190 4430 1220 4450
rect 1260 4430 1290 4450
rect 1190 4420 1290 4430
rect 1360 4450 1460 4460
rect 1360 4430 1390 4450
rect 1430 4430 1460 4450
rect 1360 4420 1460 4430
rect 1530 4450 1630 4460
rect 1530 4430 1560 4450
rect 1600 4430 1630 4450
rect 1530 4420 1630 4430
rect 1750 4450 1850 4460
rect 1750 4430 1780 4450
rect 1820 4430 1850 4450
rect 1750 4420 1850 4430
rect 1920 4450 2020 4460
rect 1920 4430 1950 4450
rect 1990 4430 2020 4450
rect 1920 4420 2020 4430
rect 2090 4450 2190 4460
rect 2090 4430 2120 4450
rect 2160 4430 2190 4450
rect 2090 4420 2190 4430
rect 2260 4450 2360 4460
rect 2260 4430 2290 4450
rect 2330 4430 2360 4450
rect 2260 4420 2360 4430
rect 2430 4450 2530 4460
rect 2430 4430 2460 4450
rect 2500 4430 2530 4450
rect 2430 4420 2530 4430
rect 2600 4450 2700 4460
rect 2600 4430 2630 4450
rect 2670 4430 2700 4450
rect 2600 4420 2700 4430
rect 2770 4450 2870 4460
rect 2770 4430 2800 4450
rect 2840 4430 2870 4450
rect 2770 4420 2870 4430
rect 2940 4450 3040 4460
rect 2940 4430 2970 4450
rect 3010 4430 3040 4450
rect 2940 4420 3040 4430
rect 3110 4450 3210 4460
rect 3110 4430 3140 4450
rect 3180 4430 3210 4450
rect 3110 4420 3210 4430
rect 3280 4450 3380 4460
rect 3280 4430 3310 4450
rect 3350 4430 3380 4450
rect 3280 4420 3380 4430
rect 0 2210 100 2220
rect 0 2190 30 2210
rect 70 2190 100 2210
rect 0 2180 100 2190
rect 170 2210 270 2220
rect 170 2190 200 2210
rect 240 2190 270 2210
rect 170 2180 270 2190
rect 340 2210 440 2220
rect 340 2190 370 2210
rect 410 2190 440 2210
rect 340 2180 440 2190
rect 510 2210 610 2220
rect 510 2190 540 2210
rect 580 2190 610 2210
rect 510 2180 610 2190
rect 680 2210 780 2220
rect 680 2190 710 2210
rect 750 2190 780 2210
rect 680 2180 780 2190
rect 850 2210 950 2220
rect 850 2190 880 2210
rect 920 2190 950 2210
rect 850 2180 950 2190
rect 1020 2210 1120 2220
rect 1020 2190 1050 2210
rect 1090 2190 1120 2210
rect 1020 2180 1120 2190
rect 1190 2210 1290 2220
rect 1190 2190 1220 2210
rect 1260 2190 1290 2210
rect 1190 2180 1290 2190
rect 1360 2210 1460 2220
rect 1360 2190 1390 2210
rect 1430 2190 1460 2210
rect 1360 2180 1460 2190
rect 1530 2210 1630 2220
rect 1530 2190 1560 2210
rect 1600 2190 1630 2210
rect 1530 2180 1630 2190
rect 1750 2210 1850 2220
rect 1750 2190 1780 2210
rect 1820 2190 1850 2210
rect 1750 2180 1850 2190
rect 1920 2210 2020 2220
rect 1920 2190 1950 2210
rect 1990 2190 2020 2210
rect 1920 2180 2020 2190
rect 2090 2210 2190 2220
rect 2090 2190 2120 2210
rect 2160 2190 2190 2210
rect 2090 2180 2190 2190
rect 2260 2210 2360 2220
rect 2260 2190 2290 2210
rect 2330 2190 2360 2210
rect 2260 2180 2360 2190
rect 2430 2210 2530 2220
rect 2430 2190 2460 2210
rect 2500 2190 2530 2210
rect 2430 2180 2530 2190
rect 2600 2210 2700 2220
rect 2600 2190 2630 2210
rect 2670 2190 2700 2210
rect 2600 2180 2700 2190
rect 2770 2210 2870 2220
rect 2770 2190 2800 2210
rect 2840 2190 2870 2210
rect 2770 2180 2870 2190
rect 2940 2210 3040 2220
rect 2940 2190 2970 2210
rect 3010 2190 3040 2210
rect 2940 2180 3040 2190
rect 3110 2210 3210 2220
rect 3110 2190 3140 2210
rect 3180 2190 3210 2210
rect 3110 2180 3210 2190
rect 3280 2210 3380 2220
rect 3280 2190 3310 2210
rect 3350 2190 3380 2210
rect 3280 2180 3380 2190
rect 0 1170 100 1180
rect 0 1150 30 1170
rect 70 1150 100 1170
rect 0 1140 100 1150
rect 170 1170 270 1180
rect 170 1150 200 1170
rect 240 1150 270 1170
rect 170 1140 270 1150
rect 340 1170 440 1180
rect 340 1150 370 1170
rect 410 1150 440 1170
rect 340 1140 440 1150
rect 510 1170 610 1180
rect 510 1150 540 1170
rect 580 1150 610 1170
rect 510 1140 610 1150
rect 680 1170 780 1180
rect 680 1150 710 1170
rect 750 1150 780 1170
rect 680 1140 780 1150
rect 850 1170 950 1180
rect 850 1150 880 1170
rect 920 1150 950 1170
rect 850 1140 950 1150
rect 1020 1170 1120 1180
rect 1020 1150 1050 1170
rect 1090 1150 1120 1170
rect 1020 1140 1120 1150
rect 1190 1170 1290 1180
rect 1190 1150 1220 1170
rect 1260 1150 1290 1170
rect 1190 1140 1290 1150
rect 1360 1170 1460 1180
rect 1360 1150 1390 1170
rect 1430 1150 1460 1170
rect 1360 1140 1460 1150
rect 1530 1170 1630 1180
rect 1530 1150 1560 1170
rect 1600 1150 1630 1170
rect 1530 1140 1630 1150
rect 1750 1170 1850 1180
rect 1750 1150 1780 1170
rect 1820 1150 1850 1170
rect 1750 1140 1850 1150
rect 1920 1170 2020 1180
rect 1920 1150 1950 1170
rect 1990 1150 2020 1170
rect 1920 1140 2020 1150
rect 2090 1170 2190 1180
rect 2090 1150 2120 1170
rect 2160 1150 2190 1170
rect 2090 1140 2190 1150
rect 2260 1170 2360 1180
rect 2260 1150 2290 1170
rect 2330 1150 2360 1170
rect 2260 1140 2360 1150
rect 2430 1170 2530 1180
rect 2430 1150 2460 1170
rect 2500 1150 2530 1170
rect 2430 1140 2530 1150
rect 2600 1170 2700 1180
rect 2600 1150 2630 1170
rect 2670 1150 2700 1170
rect 2600 1140 2700 1150
rect 2770 1170 2870 1180
rect 2770 1150 2800 1170
rect 2840 1150 2870 1170
rect 2770 1140 2870 1150
rect 2940 1170 3040 1180
rect 2940 1150 2970 1170
rect 3010 1150 3040 1170
rect 2940 1140 3040 1150
rect 3110 1170 3210 1180
rect 3110 1150 3140 1170
rect 3180 1150 3210 1170
rect 3110 1140 3210 1150
rect 3280 1170 3380 1180
rect 3280 1150 3310 1170
rect 3350 1150 3380 1170
rect 3280 1140 3380 1150
rect 0 1030 100 1040
rect 170 1030 270 1040
rect 340 1030 440 1040
rect 510 1030 610 1040
rect 680 1030 780 1040
rect 850 1030 950 1040
rect 1020 1030 1120 1040
rect 1190 1030 1290 1040
rect 1360 1030 1460 1040
rect 1530 1030 1630 1040
rect 1750 1030 1850 1040
rect 1920 1030 2020 1040
rect 2090 1030 2190 1040
rect 2260 1030 2360 1040
rect 2430 1030 2530 1040
rect 2600 1030 2700 1040
rect 2770 1030 2870 1040
rect 2940 1030 3040 1040
rect 3110 1030 3210 1040
rect 3280 1030 3380 1040
rect 0 1010 30 1030
rect 70 1010 200 1030
rect 240 1010 370 1030
rect 410 1010 540 1030
rect 580 1010 710 1030
rect 750 1010 880 1030
rect 920 1010 1050 1030
rect 1090 1010 1220 1030
rect 1260 1010 1390 1030
rect 1430 1010 1560 1030
rect 1600 1010 1780 1030
rect 1820 1010 1950 1030
rect 1990 1010 2120 1030
rect 2160 1010 2290 1030
rect 2330 1010 2460 1030
rect 2500 1010 2630 1030
rect 2670 1010 2800 1030
rect 2840 1010 2970 1030
rect 3010 1010 3140 1030
rect 3180 1010 3310 1030
rect 3350 1010 3380 1030
rect 0 1000 100 1010
rect 170 1000 270 1010
rect 340 1000 440 1010
rect 510 1000 610 1010
rect 680 1000 780 1010
rect 850 1000 950 1010
rect 1020 1000 1120 1010
rect 1190 1000 1290 1010
rect 1360 1000 1460 1010
rect 1530 1000 1630 1010
rect 1750 1000 1850 1010
rect 1920 1000 2020 1010
rect 2090 1000 2190 1010
rect 2260 1000 2360 1010
rect 2430 1000 2530 1010
rect 2600 1000 2700 1010
rect 2770 1000 2870 1010
rect 2940 1000 3040 1010
rect 3110 1000 3210 1010
rect 3280 1000 3380 1010
rect 0 890 100 900
rect 0 870 30 890
rect 70 870 100 890
rect 0 860 100 870
rect 170 890 270 900
rect 170 870 200 890
rect 240 870 270 890
rect 170 860 270 870
rect 340 890 440 900
rect 340 870 370 890
rect 410 870 440 890
rect 340 860 440 870
rect 510 890 610 900
rect 510 870 540 890
rect 580 870 610 890
rect 510 860 610 870
rect 680 890 780 900
rect 680 870 710 890
rect 750 870 780 890
rect 680 860 780 870
rect 850 890 950 900
rect 850 870 880 890
rect 920 870 950 890
rect 850 860 950 870
rect 1020 890 1120 900
rect 1020 870 1050 890
rect 1090 870 1120 890
rect 1020 860 1120 870
rect 1190 890 1290 900
rect 1190 870 1220 890
rect 1260 870 1290 890
rect 1190 860 1290 870
rect 1360 890 1460 900
rect 1360 870 1390 890
rect 1430 870 1460 890
rect 1360 860 1460 870
rect 1530 890 1630 900
rect 1530 870 1560 890
rect 1600 870 1630 890
rect 1530 860 1630 870
rect 1750 890 1850 900
rect 1750 870 1780 890
rect 1820 870 1850 890
rect 1750 860 1850 870
rect 1920 890 2020 900
rect 1920 870 1950 890
rect 1990 870 2020 890
rect 1920 860 2020 870
rect 2090 890 2190 900
rect 2090 870 2120 890
rect 2160 870 2190 890
rect 2090 860 2190 870
rect 2260 890 2360 900
rect 2260 870 2290 890
rect 2330 870 2360 890
rect 2260 860 2360 870
rect 2430 890 2530 900
rect 2430 870 2460 890
rect 2500 870 2530 890
rect 2430 860 2530 870
rect 2600 890 2700 900
rect 2600 870 2630 890
rect 2670 870 2700 890
rect 2600 860 2700 870
rect 2770 890 2870 900
rect 2770 870 2800 890
rect 2840 870 2870 890
rect 2770 860 2870 870
rect 2940 890 3040 900
rect 2940 870 2970 890
rect 3010 870 3040 890
rect 2940 860 3040 870
rect 3110 890 3210 900
rect 3110 870 3140 890
rect 3180 870 3210 890
rect 3110 860 3210 870
rect 3280 890 3380 900
rect 3280 870 3310 890
rect 3350 870 3380 890
rect 3280 860 3380 870
<< ndiffc >>
rect -200 5610 -160 5630
rect 3540 5610 3580 5630
rect -200 5070 -160 5090
rect -220 4530 -180 4550
rect 3540 5070 3580 5090
rect 3560 4530 3600 4550
rect -190 3820 -170 3860
rect -50 3820 -30 3860
rect 90 3820 110 3860
rect 230 3820 250 3860
rect 370 3820 390 3860
rect 510 3820 530 3860
rect 650 3820 670 3860
rect 790 3820 810 3860
rect 930 3820 950 3860
rect 1070 3820 1090 3860
rect 1210 3820 1230 3860
rect 1560 4310 1580 4330
rect 1800 4310 1820 4330
rect 1350 3820 1370 3860
rect 1560 3830 1580 3850
rect 1800 3830 1820 3850
rect 2010 3820 2030 3860
rect -190 2780 -170 2820
rect -50 2780 -30 2820
rect 90 2780 110 2820
rect 230 2780 250 2820
rect 370 2780 390 2820
rect 510 2780 530 2820
rect 650 2780 670 2820
rect 790 2780 810 2820
rect 930 2780 950 2820
rect 1070 2780 1090 2820
rect 1210 2780 1230 2820
rect 1560 3310 1580 3330
rect 1800 3310 1820 3330
rect 2150 3820 2170 3860
rect 2290 3820 2310 3860
rect 2430 3820 2450 3860
rect 2570 3820 2590 3860
rect 2710 3820 2730 3860
rect 2850 3820 2870 3860
rect 2990 3820 3010 3860
rect 3130 3820 3150 3860
rect 3270 3820 3290 3860
rect 3410 3820 3430 3860
rect 3550 3820 3570 3860
rect 1350 2780 1370 2820
rect 1560 2790 1580 2810
rect 1800 2790 1820 2810
rect 2010 2780 2030 2820
rect 1560 2310 1580 2330
rect 1800 2310 1820 2330
rect 2150 2780 2170 2820
rect 2290 2780 2310 2820
rect 2430 2780 2450 2820
rect 2570 2780 2590 2820
rect 2710 2780 2730 2820
rect 2850 2780 2870 2820
rect 2990 2780 3010 2820
rect 3130 2780 3150 2820
rect 3270 2780 3290 2820
rect 3410 2780 3430 2820
rect 3550 2780 3570 2820
rect -220 2090 -180 2110
rect -200 1550 -160 1570
rect 3560 2090 3600 2110
rect 3540 1550 3580 1570
rect -200 1010 -160 1030
rect 3540 1010 3580 1030
<< pdiffc >>
rect 30 5750 70 5770
rect 200 5750 240 5770
rect 370 5750 410 5770
rect 540 5750 580 5770
rect 710 5750 750 5770
rect 880 5750 920 5770
rect 1050 5750 1090 5770
rect 1220 5750 1260 5770
rect 1390 5750 1430 5770
rect 1560 5750 1600 5770
rect 1780 5750 1820 5770
rect 1950 5750 1990 5770
rect 2120 5750 2160 5770
rect 2290 5750 2330 5770
rect 2460 5750 2500 5770
rect 2630 5750 2670 5770
rect 2800 5750 2840 5770
rect 2970 5750 3010 5770
rect 3140 5750 3180 5770
rect 3310 5750 3350 5770
rect 30 5610 70 5630
rect 200 5610 240 5630
rect 370 5610 410 5630
rect 540 5610 580 5630
rect 710 5610 750 5630
rect 880 5610 920 5630
rect 1050 5610 1090 5630
rect 1220 5610 1260 5630
rect 1390 5610 1430 5630
rect 1560 5610 1600 5630
rect 1780 5610 1820 5630
rect 1950 5610 1990 5630
rect 2120 5610 2160 5630
rect 2290 5610 2330 5630
rect 2460 5610 2500 5630
rect 2630 5610 2670 5630
rect 2800 5610 2840 5630
rect 2970 5610 3010 5630
rect 3140 5610 3180 5630
rect 3310 5610 3350 5630
rect 30 5470 70 5490
rect 200 5470 240 5490
rect 370 5470 410 5490
rect 540 5470 580 5490
rect 710 5470 750 5490
rect 880 5470 920 5490
rect 1050 5470 1090 5490
rect 1220 5470 1260 5490
rect 1390 5470 1430 5490
rect 1560 5470 1600 5490
rect 1780 5470 1820 5490
rect 1950 5470 1990 5490
rect 2120 5470 2160 5490
rect 2290 5470 2330 5490
rect 2460 5470 2500 5490
rect 2630 5470 2670 5490
rect 2800 5470 2840 5490
rect 2970 5470 3010 5490
rect 3140 5470 3180 5490
rect 3310 5470 3350 5490
rect 30 4430 70 4450
rect 200 4430 240 4450
rect 370 4430 410 4450
rect 540 4430 580 4450
rect 710 4430 750 4450
rect 880 4430 920 4450
rect 1050 4430 1090 4450
rect 1220 4430 1260 4450
rect 1390 4430 1430 4450
rect 1560 4430 1600 4450
rect 1780 4430 1820 4450
rect 1950 4430 1990 4450
rect 2120 4430 2160 4450
rect 2290 4430 2330 4450
rect 2460 4430 2500 4450
rect 2630 4430 2670 4450
rect 2800 4430 2840 4450
rect 2970 4430 3010 4450
rect 3140 4430 3180 4450
rect 3310 4430 3350 4450
rect 30 2190 70 2210
rect 200 2190 240 2210
rect 370 2190 410 2210
rect 540 2190 580 2210
rect 710 2190 750 2210
rect 880 2190 920 2210
rect 1050 2190 1090 2210
rect 1220 2190 1260 2210
rect 1390 2190 1430 2210
rect 1560 2190 1600 2210
rect 1780 2190 1820 2210
rect 1950 2190 1990 2210
rect 2120 2190 2160 2210
rect 2290 2190 2330 2210
rect 2460 2190 2500 2210
rect 2630 2190 2670 2210
rect 2800 2190 2840 2210
rect 2970 2190 3010 2210
rect 3140 2190 3180 2210
rect 3310 2190 3350 2210
rect 30 1150 70 1170
rect 200 1150 240 1170
rect 370 1150 410 1170
rect 540 1150 580 1170
rect 710 1150 750 1170
rect 880 1150 920 1170
rect 1050 1150 1090 1170
rect 1220 1150 1260 1170
rect 1390 1150 1430 1170
rect 1560 1150 1600 1170
rect 1780 1150 1820 1170
rect 1950 1150 1990 1170
rect 2120 1150 2160 1170
rect 2290 1150 2330 1170
rect 2460 1150 2500 1170
rect 2630 1150 2670 1170
rect 2800 1150 2840 1170
rect 2970 1150 3010 1170
rect 3140 1150 3180 1170
rect 3310 1150 3350 1170
rect 30 1010 70 1030
rect 200 1010 240 1030
rect 370 1010 410 1030
rect 540 1010 580 1030
rect 710 1010 750 1030
rect 880 1010 920 1030
rect 1050 1010 1090 1030
rect 1220 1010 1260 1030
rect 1390 1010 1430 1030
rect 1560 1010 1600 1030
rect 1780 1010 1820 1030
rect 1950 1010 1990 1030
rect 2120 1010 2160 1030
rect 2290 1010 2330 1030
rect 2460 1010 2500 1030
rect 2630 1010 2670 1030
rect 2800 1010 2840 1030
rect 2970 1010 3010 1030
rect 3140 1010 3180 1030
rect 3310 1010 3350 1030
rect 30 870 70 890
rect 200 870 240 890
rect 370 870 410 890
rect 540 870 580 890
rect 710 870 750 890
rect 880 870 920 890
rect 1050 870 1090 890
rect 1220 870 1260 890
rect 1390 870 1430 890
rect 1560 870 1600 890
rect 1780 870 1820 890
rect 1950 870 1990 890
rect 2120 870 2160 890
rect 2290 870 2330 890
rect 2460 870 2500 890
rect 2630 870 2670 890
rect 2800 870 2840 890
rect 2970 870 3010 890
rect 3140 870 3180 890
rect 3310 870 3350 890
<< psubdiff >>
rect -240 4310 -200 4320
rect -240 4270 -230 4310
rect -210 4270 -200 4310
rect -240 4260 -200 4270
rect 1440 3330 1500 3350
rect 1440 3310 1460 3330
rect 1480 3310 1500 3330
rect -240 2370 -200 2380
rect -240 2330 -230 2370
rect -210 2330 -200 2370
rect -240 2320 -200 2330
rect 1440 3290 1500 3310
rect 1880 3330 1940 3350
rect 3580 4310 3620 4320
rect 3580 4270 3590 4310
rect 3610 4270 3620 4310
rect 3580 4260 3620 4270
rect 1880 3310 1900 3330
rect 1920 3310 1940 3330
rect 1880 3290 1940 3310
rect 3580 2370 3620 2380
rect 3580 2330 3590 2370
rect 3610 2330 3620 2370
rect 3580 2320 3620 2330
<< nsubdiff >>
rect 0 5790 30 5810
rect 70 5790 100 5810
rect 0 5780 100 5790
rect 170 5790 200 5810
rect 240 5790 270 5810
rect 170 5780 270 5790
rect 340 5790 370 5810
rect 410 5790 440 5810
rect 340 5780 440 5790
rect 510 5790 540 5810
rect 580 5790 610 5810
rect 510 5780 610 5790
rect 680 5790 710 5810
rect 750 5790 780 5810
rect 680 5780 780 5790
rect 850 5790 880 5810
rect 920 5790 950 5810
rect 850 5780 950 5790
rect 1020 5790 1050 5810
rect 1090 5790 1120 5810
rect 1020 5780 1120 5790
rect 1190 5790 1220 5810
rect 1260 5790 1290 5810
rect 1190 5780 1290 5790
rect 1360 5790 1390 5810
rect 1430 5790 1460 5810
rect 1360 5780 1460 5790
rect 1530 5790 1560 5810
rect 1600 5790 1630 5810
rect 1530 5780 1630 5790
rect 1750 5790 1780 5810
rect 1820 5790 1850 5810
rect 1750 5780 1850 5790
rect 1920 5790 1950 5810
rect 1990 5790 2020 5810
rect 1920 5780 2020 5790
rect 2090 5790 2120 5810
rect 2160 5790 2190 5810
rect 2090 5780 2190 5790
rect 2260 5790 2290 5810
rect 2330 5790 2360 5810
rect 2260 5780 2360 5790
rect 2430 5790 2460 5810
rect 2500 5790 2530 5810
rect 2430 5780 2530 5790
rect 2600 5790 2630 5810
rect 2670 5790 2700 5810
rect 2600 5780 2700 5790
rect 2770 5790 2800 5810
rect 2840 5790 2870 5810
rect 2770 5780 2870 5790
rect 2940 5790 2970 5810
rect 3010 5790 3040 5810
rect 2940 5780 3040 5790
rect 3110 5790 3140 5810
rect 3180 5790 3210 5810
rect 3110 5780 3210 5790
rect 3280 5790 3310 5810
rect 3350 5790 3380 5810
rect 3280 5780 3380 5790
rect 0 850 100 860
rect 0 830 30 850
rect 70 830 100 850
rect 170 850 270 860
rect 170 830 200 850
rect 240 830 270 850
rect 340 850 440 860
rect 340 830 370 850
rect 410 830 440 850
rect 510 850 610 860
rect 510 830 540 850
rect 580 830 610 850
rect 680 850 780 860
rect 680 830 710 850
rect 750 830 780 850
rect 850 850 950 860
rect 850 830 880 850
rect 920 830 950 850
rect 1020 850 1120 860
rect 1020 830 1050 850
rect 1090 830 1120 850
rect 1190 850 1290 860
rect 1190 830 1220 850
rect 1260 830 1290 850
rect 1360 850 1460 860
rect 1360 830 1390 850
rect 1430 830 1460 850
rect 1530 850 1630 860
rect 1530 830 1560 850
rect 1600 830 1630 850
rect 1750 850 1850 860
rect 1750 830 1780 850
rect 1820 830 1850 850
rect 1920 850 2020 860
rect 1920 830 1950 850
rect 1990 830 2020 850
rect 2090 850 2190 860
rect 2090 830 2120 850
rect 2160 830 2190 850
rect 2260 850 2360 860
rect 2260 830 2290 850
rect 2330 830 2360 850
rect 2430 850 2530 860
rect 2430 830 2460 850
rect 2500 830 2530 850
rect 2600 850 2700 860
rect 2600 830 2630 850
rect 2670 830 2700 850
rect 2770 850 2870 860
rect 2770 830 2800 850
rect 2840 830 2870 850
rect 2940 850 3040 860
rect 2940 830 2970 850
rect 3010 830 3040 850
rect 3110 850 3210 860
rect 3110 830 3140 850
rect 3180 830 3210 850
rect 3280 850 3380 860
rect 3280 830 3310 850
rect 3350 830 3380 850
<< psubdiffcont >>
rect -230 4270 -210 4310
rect 1460 3310 1480 3330
rect -230 2330 -210 2370
rect 3590 4270 3610 4310
rect 1900 3310 1920 3330
rect 3590 2330 3610 2370
<< nsubdiffcont >>
rect 30 5790 70 5810
rect 200 5790 240 5810
rect 370 5790 410 5810
rect 540 5790 580 5810
rect 710 5790 750 5810
rect 880 5790 920 5810
rect 1050 5790 1090 5810
rect 1220 5790 1260 5810
rect 1390 5790 1430 5810
rect 1560 5790 1600 5810
rect 1780 5790 1820 5810
rect 1950 5790 1990 5810
rect 2120 5790 2160 5810
rect 2290 5790 2330 5810
rect 2460 5790 2500 5810
rect 2630 5790 2670 5810
rect 2800 5790 2840 5810
rect 2970 5790 3010 5810
rect 3140 5790 3180 5810
rect 3310 5790 3350 5810
rect 30 830 70 850
rect 200 830 240 850
rect 370 830 410 850
rect 540 830 580 850
rect 710 830 750 850
rect 880 830 920 850
rect 1050 830 1090 850
rect 1220 830 1260 850
rect 1390 830 1430 850
rect 1560 830 1600 850
rect 1780 830 1820 850
rect 1950 830 1990 850
rect 2120 830 2160 850
rect 2290 830 2330 850
rect 2460 830 2500 850
rect 2630 830 2670 850
rect 2800 830 2840 850
rect 2970 830 3010 850
rect 3140 830 3180 850
rect 3310 830 3350 850
<< poly >>
rect -60 5790 -20 5800
rect -60 5770 -50 5790
rect -30 5770 -20 5790
rect -60 5740 -20 5770
rect 3400 5790 3440 5800
rect 3400 5770 3410 5790
rect 3430 5770 3440 5790
rect 3400 5740 3440 5770
rect -310 5690 -270 5700
rect -310 5670 -300 5690
rect -280 5670 -270 5690
rect -310 5660 -270 5670
rect -310 5600 -290 5660
rect -60 5640 0 5740
rect 100 5710 120 5740
rect 150 5710 170 5740
rect 100 5670 170 5710
rect 100 5640 120 5670
rect 150 5640 170 5670
rect 270 5710 290 5740
rect 320 5710 340 5740
rect 270 5670 340 5710
rect 270 5640 290 5670
rect 320 5640 340 5670
rect 440 5710 460 5740
rect 490 5710 510 5740
rect 440 5670 510 5710
rect 440 5640 460 5670
rect 490 5640 510 5670
rect 610 5710 630 5740
rect 660 5710 680 5740
rect 610 5670 680 5710
rect 610 5640 630 5670
rect 660 5640 680 5670
rect 780 5710 800 5740
rect 830 5710 850 5740
rect 780 5670 850 5710
rect 780 5640 800 5670
rect 830 5640 850 5670
rect 950 5710 970 5740
rect 1000 5710 1020 5740
rect 950 5670 1020 5710
rect 950 5640 970 5670
rect 1000 5640 1020 5670
rect 1120 5710 1140 5740
rect 1170 5710 1190 5740
rect 1120 5670 1190 5710
rect 1120 5640 1140 5670
rect 1170 5640 1190 5670
rect 1290 5710 1310 5740
rect 1340 5710 1360 5740
rect 1290 5670 1360 5710
rect 1290 5640 1310 5670
rect 1340 5640 1360 5670
rect 1460 5710 1480 5740
rect 1510 5710 1530 5740
rect 1460 5670 1530 5710
rect 1460 5640 1480 5670
rect 1510 5640 1530 5670
rect 1630 5710 1650 5740
rect 1730 5710 1750 5740
rect 1630 5670 1750 5710
rect 1630 5640 1650 5670
rect 1730 5640 1750 5670
rect 1850 5710 1870 5740
rect 1900 5710 1920 5740
rect 1850 5670 1920 5710
rect 1850 5640 1870 5670
rect 1900 5640 1920 5670
rect 2020 5710 2040 5740
rect 2070 5710 2090 5740
rect 2020 5670 2090 5710
rect 2020 5640 2040 5670
rect 2070 5640 2090 5670
rect 2190 5710 2210 5740
rect 2240 5710 2260 5740
rect 2190 5670 2260 5710
rect 2190 5640 2210 5670
rect 2240 5640 2260 5670
rect 2360 5710 2380 5740
rect 2410 5710 2430 5740
rect 2360 5670 2430 5710
rect 2360 5640 2380 5670
rect 2410 5640 2430 5670
rect 2530 5710 2550 5740
rect 2580 5710 2600 5740
rect 2530 5670 2600 5710
rect 2530 5640 2550 5670
rect 2580 5640 2600 5670
rect 2700 5710 2720 5740
rect 2750 5710 2770 5740
rect 2700 5670 2770 5710
rect 2700 5640 2720 5670
rect 2750 5640 2770 5670
rect 2870 5710 2890 5740
rect 2920 5710 2940 5740
rect 2870 5670 2940 5710
rect 2870 5640 2890 5670
rect 2920 5640 2940 5670
rect 3040 5710 3060 5740
rect 3090 5710 3110 5740
rect 3040 5670 3110 5710
rect 3040 5640 3060 5670
rect 3090 5640 3110 5670
rect 3210 5710 3230 5740
rect 3260 5710 3280 5740
rect 3210 5670 3280 5710
rect 3210 5640 3230 5670
rect 3260 5640 3280 5670
rect 3380 5640 3440 5740
rect 3650 5690 3690 5700
rect 3650 5670 3660 5690
rect 3680 5670 3690 5690
rect 3650 5660 3690 5670
rect 3670 5600 3690 5660
rect -310 5100 -280 5600
rect -80 5100 -60 5600
rect -20 5500 0 5600
rect 100 5570 120 5600
rect 150 5570 170 5600
rect 100 5530 170 5570
rect 100 5500 120 5530
rect 150 5500 170 5530
rect 270 5570 290 5600
rect 320 5570 340 5600
rect 270 5530 340 5570
rect 270 5500 290 5530
rect 320 5500 340 5530
rect 440 5570 460 5600
rect 490 5570 510 5600
rect 440 5530 510 5570
rect 440 5500 460 5530
rect 490 5500 510 5530
rect 610 5570 630 5600
rect 660 5570 680 5600
rect 610 5530 680 5570
rect 610 5500 630 5530
rect 660 5500 680 5530
rect 780 5570 800 5600
rect 830 5570 850 5600
rect 780 5530 850 5570
rect 780 5500 800 5530
rect 830 5500 850 5530
rect 950 5570 970 5600
rect 1000 5570 1020 5600
rect 950 5530 1020 5570
rect 950 5500 970 5530
rect 1000 5500 1020 5530
rect 1120 5570 1140 5600
rect 1170 5570 1190 5600
rect 1120 5530 1190 5570
rect 1120 5500 1140 5530
rect 1170 5500 1190 5530
rect 1290 5570 1310 5600
rect 1340 5570 1360 5600
rect 1290 5530 1360 5570
rect 1290 5500 1310 5530
rect 1340 5500 1360 5530
rect 1460 5570 1480 5600
rect 1510 5570 1530 5600
rect 1460 5530 1530 5570
rect 1460 5500 1480 5530
rect 1510 5500 1530 5530
rect 1630 5570 1650 5600
rect 1730 5570 1750 5600
rect 1630 5530 1750 5570
rect 1630 5500 1650 5530
rect -300 4560 -280 5060
rect -80 4560 -50 5060
rect -70 4500 -50 4560
rect -90 4490 -50 4500
rect -90 4470 -80 4490
rect -60 4470 -50 4490
rect -90 4460 -50 4470
rect -20 4460 0 5460
rect 100 5430 120 5460
rect 150 5430 170 5460
rect 100 5390 170 5430
rect 100 5330 120 5390
rect 150 5330 170 5390
rect 100 5290 170 5330
rect 100 5230 120 5290
rect 150 5230 170 5290
rect 100 5190 170 5230
rect 100 5130 120 5190
rect 150 5130 170 5190
rect 100 5090 170 5130
rect 100 5030 120 5090
rect 150 5030 170 5090
rect 100 4990 170 5030
rect 100 4930 120 4990
rect 150 4930 170 4990
rect 100 4890 170 4930
rect 100 4830 120 4890
rect 150 4830 170 4890
rect 100 4790 170 4830
rect 100 4730 120 4790
rect 150 4730 170 4790
rect 100 4690 170 4730
rect 100 4630 120 4690
rect 150 4630 170 4690
rect 100 4590 170 4630
rect 100 4530 120 4590
rect 150 4530 170 4590
rect 100 4490 170 4530
rect 100 4460 120 4490
rect 150 4460 170 4490
rect 270 5430 290 5460
rect 320 5430 340 5460
rect 270 5390 340 5430
rect 270 5330 290 5390
rect 320 5330 340 5390
rect 270 5290 340 5330
rect 270 5230 290 5290
rect 320 5230 340 5290
rect 270 5190 340 5230
rect 270 5130 290 5190
rect 320 5130 340 5190
rect 270 5090 340 5130
rect 270 5030 290 5090
rect 320 5030 340 5090
rect 270 4990 340 5030
rect 270 4930 290 4990
rect 320 4930 340 4990
rect 270 4890 340 4930
rect 270 4830 290 4890
rect 320 4830 340 4890
rect 270 4790 340 4830
rect 270 4730 290 4790
rect 320 4730 340 4790
rect 270 4690 340 4730
rect 270 4630 290 4690
rect 320 4630 340 4690
rect 270 4590 340 4630
rect 270 4530 290 4590
rect 320 4530 340 4590
rect 270 4490 340 4530
rect 270 4460 290 4490
rect 320 4460 340 4490
rect 440 5430 460 5460
rect 490 5430 510 5460
rect 440 5390 510 5430
rect 440 5330 460 5390
rect 490 5330 510 5390
rect 440 5290 510 5330
rect 440 5230 460 5290
rect 490 5230 510 5290
rect 440 5190 510 5230
rect 440 5130 460 5190
rect 490 5130 510 5190
rect 440 5090 510 5130
rect 440 5030 460 5090
rect 490 5030 510 5090
rect 440 4990 510 5030
rect 440 4930 460 4990
rect 490 4930 510 4990
rect 440 4890 510 4930
rect 440 4830 460 4890
rect 490 4830 510 4890
rect 440 4790 510 4830
rect 440 4730 460 4790
rect 490 4730 510 4790
rect 440 4690 510 4730
rect 440 4630 460 4690
rect 490 4630 510 4690
rect 440 4590 510 4630
rect 440 4530 460 4590
rect 490 4530 510 4590
rect 440 4490 510 4530
rect 440 4460 460 4490
rect 490 4460 510 4490
rect 610 5430 630 5460
rect 660 5430 680 5460
rect 610 5390 680 5430
rect 610 5330 630 5390
rect 660 5330 680 5390
rect 610 5290 680 5330
rect 610 5230 630 5290
rect 660 5230 680 5290
rect 610 5190 680 5230
rect 610 5130 630 5190
rect 660 5130 680 5190
rect 610 5090 680 5130
rect 610 5030 630 5090
rect 660 5030 680 5090
rect 610 4990 680 5030
rect 610 4930 630 4990
rect 660 4930 680 4990
rect 610 4890 680 4930
rect 610 4830 630 4890
rect 660 4830 680 4890
rect 610 4790 680 4830
rect 610 4730 630 4790
rect 660 4730 680 4790
rect 610 4690 680 4730
rect 610 4630 630 4690
rect 660 4630 680 4690
rect 610 4590 680 4630
rect 610 4530 630 4590
rect 660 4530 680 4590
rect 610 4490 680 4530
rect 610 4460 630 4490
rect 660 4460 680 4490
rect 780 5430 800 5460
rect 830 5430 850 5460
rect 780 5390 850 5430
rect 780 5330 800 5390
rect 830 5330 850 5390
rect 780 5290 850 5330
rect 780 5230 800 5290
rect 830 5230 850 5290
rect 780 5190 850 5230
rect 780 5130 800 5190
rect 830 5130 850 5190
rect 780 5090 850 5130
rect 780 5030 800 5090
rect 830 5030 850 5090
rect 780 4990 850 5030
rect 780 4930 800 4990
rect 830 4930 850 4990
rect 780 4890 850 4930
rect 780 4830 800 4890
rect 830 4830 850 4890
rect 780 4790 850 4830
rect 780 4730 800 4790
rect 830 4730 850 4790
rect 780 4690 850 4730
rect 780 4630 800 4690
rect 830 4630 850 4690
rect 780 4590 850 4630
rect 780 4530 800 4590
rect 830 4530 850 4590
rect 780 4490 850 4530
rect 780 4460 800 4490
rect 830 4460 850 4490
rect 950 5430 970 5460
rect 1000 5430 1020 5460
rect 950 5390 1020 5430
rect 950 5330 970 5390
rect 1000 5330 1020 5390
rect 950 5290 1020 5330
rect 950 5230 970 5290
rect 1000 5230 1020 5290
rect 950 5190 1020 5230
rect 950 5130 970 5190
rect 1000 5130 1020 5190
rect 950 5090 1020 5130
rect 950 5030 970 5090
rect 1000 5030 1020 5090
rect 950 4990 1020 5030
rect 950 4930 970 4990
rect 1000 4930 1020 4990
rect 950 4890 1020 4930
rect 950 4830 970 4890
rect 1000 4830 1020 4890
rect 950 4790 1020 4830
rect 950 4730 970 4790
rect 1000 4730 1020 4790
rect 950 4690 1020 4730
rect 950 4630 970 4690
rect 1000 4630 1020 4690
rect 950 4590 1020 4630
rect 950 4530 970 4590
rect 1000 4530 1020 4590
rect 950 4490 1020 4530
rect 950 4460 970 4490
rect 1000 4460 1020 4490
rect 1120 5430 1140 5460
rect 1170 5430 1190 5460
rect 1120 5390 1190 5430
rect 1120 5330 1140 5390
rect 1170 5330 1190 5390
rect 1120 5290 1190 5330
rect 1120 5230 1140 5290
rect 1170 5230 1190 5290
rect 1120 5190 1190 5230
rect 1120 5130 1140 5190
rect 1170 5130 1190 5190
rect 1120 5090 1190 5130
rect 1120 5030 1140 5090
rect 1170 5030 1190 5090
rect 1120 4990 1190 5030
rect 1120 4930 1140 4990
rect 1170 4930 1190 4990
rect 1120 4890 1190 4930
rect 1120 4830 1140 4890
rect 1170 4830 1190 4890
rect 1120 4790 1190 4830
rect 1120 4730 1140 4790
rect 1170 4730 1190 4790
rect 1120 4690 1190 4730
rect 1120 4630 1140 4690
rect 1170 4630 1190 4690
rect 1120 4590 1190 4630
rect 1120 4530 1140 4590
rect 1170 4530 1190 4590
rect 1120 4490 1190 4530
rect 1120 4460 1140 4490
rect 1170 4460 1190 4490
rect 1290 5430 1310 5460
rect 1340 5430 1360 5460
rect 1290 5390 1360 5430
rect 1290 5330 1310 5390
rect 1340 5330 1360 5390
rect 1290 5290 1360 5330
rect 1290 5230 1310 5290
rect 1340 5230 1360 5290
rect 1290 5190 1360 5230
rect 1290 5130 1310 5190
rect 1340 5130 1360 5190
rect 1290 5090 1360 5130
rect 1290 5030 1310 5090
rect 1340 5030 1360 5090
rect 1290 4990 1360 5030
rect 1290 4930 1310 4990
rect 1340 4930 1360 4990
rect 1290 4890 1360 4930
rect 1290 4830 1310 4890
rect 1340 4830 1360 4890
rect 1290 4790 1360 4830
rect 1290 4730 1310 4790
rect 1340 4730 1360 4790
rect 1290 4690 1360 4730
rect 1290 4630 1310 4690
rect 1340 4630 1360 4690
rect 1290 4590 1360 4630
rect 1290 4530 1310 4590
rect 1340 4530 1360 4590
rect 1290 4490 1360 4530
rect 1290 4460 1310 4490
rect 1340 4460 1360 4490
rect 1460 5430 1480 5460
rect 1510 5430 1530 5460
rect 1460 5390 1530 5430
rect 1460 5330 1480 5390
rect 1510 5330 1530 5390
rect 1460 5290 1530 5330
rect 1460 5230 1480 5290
rect 1510 5230 1530 5290
rect 1460 5190 1530 5230
rect 1460 5130 1480 5190
rect 1510 5130 1530 5190
rect 1460 5090 1530 5130
rect 1460 5030 1480 5090
rect 1510 5030 1530 5090
rect 1460 4990 1530 5030
rect 1460 4930 1480 4990
rect 1510 4930 1530 4990
rect 1460 4890 1530 4930
rect 1460 4830 1480 4890
rect 1510 4830 1530 4890
rect 1460 4790 1530 4830
rect 1460 4730 1480 4790
rect 1510 4730 1530 4790
rect 1460 4690 1530 4730
rect 1460 4630 1480 4690
rect 1510 4630 1530 4690
rect 1460 4590 1530 4630
rect 1460 4530 1480 4590
rect 1510 4530 1530 4590
rect 1460 4490 1530 4530
rect 1460 4460 1480 4490
rect 1510 4460 1530 4490
rect 1630 5430 1650 5460
rect 1680 5430 1700 5530
rect 1730 5500 1750 5530
rect 1850 5570 1870 5600
rect 1900 5570 1920 5600
rect 1850 5530 1920 5570
rect 1850 5500 1870 5530
rect 1900 5500 1920 5530
rect 2020 5570 2040 5600
rect 2070 5570 2090 5600
rect 2020 5530 2090 5570
rect 2020 5500 2040 5530
rect 2070 5500 2090 5530
rect 2190 5570 2210 5600
rect 2240 5570 2260 5600
rect 2190 5530 2260 5570
rect 2190 5500 2210 5530
rect 2240 5500 2260 5530
rect 2360 5570 2380 5600
rect 2410 5570 2430 5600
rect 2360 5530 2430 5570
rect 2360 5500 2380 5530
rect 2410 5500 2430 5530
rect 2530 5570 2550 5600
rect 2580 5570 2600 5600
rect 2530 5530 2600 5570
rect 2530 5500 2550 5530
rect 2580 5500 2600 5530
rect 2700 5570 2720 5600
rect 2750 5570 2770 5600
rect 2700 5530 2770 5570
rect 2700 5500 2720 5530
rect 2750 5500 2770 5530
rect 2870 5570 2890 5600
rect 2920 5570 2940 5600
rect 2870 5530 2940 5570
rect 2870 5500 2890 5530
rect 2920 5500 2940 5530
rect 3040 5570 3060 5600
rect 3090 5570 3110 5600
rect 3040 5530 3110 5570
rect 3040 5500 3060 5530
rect 3090 5500 3110 5530
rect 3210 5570 3230 5600
rect 3260 5570 3280 5600
rect 3210 5530 3280 5570
rect 3210 5500 3230 5530
rect 3260 5500 3280 5530
rect 3380 5500 3400 5600
rect 1730 5430 1750 5460
rect 1630 5390 1750 5430
rect 1630 5330 1650 5390
rect 1680 5330 1700 5390
rect 1730 5330 1750 5390
rect 1630 5290 1750 5330
rect 1630 5230 1650 5290
rect 1680 5230 1700 5290
rect 1730 5230 1750 5290
rect 1630 5190 1750 5230
rect 1630 5130 1650 5190
rect 1680 5130 1700 5190
rect 1730 5130 1750 5190
rect 1630 5090 1750 5130
rect 1630 5030 1650 5090
rect 1680 5030 1700 5090
rect 1730 5030 1750 5090
rect 1630 4990 1750 5030
rect 1630 4930 1650 4990
rect 1680 4930 1700 4990
rect 1730 4930 1750 4990
rect 1630 4890 1750 4930
rect 1630 4830 1650 4890
rect 1680 4830 1700 4890
rect 1730 4830 1750 4890
rect 1630 4790 1750 4830
rect 1630 4730 1650 4790
rect 1680 4730 1700 4790
rect 1730 4730 1750 4790
rect 1630 4690 1750 4730
rect 1630 4630 1650 4690
rect 1680 4630 1700 4690
rect 1730 4630 1750 4690
rect 1630 4590 1750 4630
rect 1630 4530 1650 4590
rect 1680 4530 1700 4590
rect 1730 4530 1750 4590
rect 1630 4490 1750 4530
rect 1630 4460 1650 4490
rect 1680 4400 1700 4490
rect 1730 4460 1750 4490
rect 1850 5430 1870 5460
rect 1900 5430 1920 5460
rect 1850 5390 1920 5430
rect 1850 5330 1870 5390
rect 1900 5330 1920 5390
rect 1850 5290 1920 5330
rect 1850 5230 1870 5290
rect 1900 5230 1920 5290
rect 1850 5190 1920 5230
rect 1850 5130 1870 5190
rect 1900 5130 1920 5190
rect 1850 5090 1920 5130
rect 1850 5030 1870 5090
rect 1900 5030 1920 5090
rect 1850 4990 1920 5030
rect 1850 4930 1870 4990
rect 1900 4930 1920 4990
rect 1850 4890 1920 4930
rect 1850 4830 1870 4890
rect 1900 4830 1920 4890
rect 1850 4790 1920 4830
rect 1850 4730 1870 4790
rect 1900 4730 1920 4790
rect 1850 4690 1920 4730
rect 1850 4630 1870 4690
rect 1900 4630 1920 4690
rect 1850 4590 1920 4630
rect 1850 4530 1870 4590
rect 1900 4530 1920 4590
rect 1850 4490 1920 4530
rect 1850 4460 1870 4490
rect 1900 4460 1920 4490
rect 2020 5430 2040 5460
rect 2070 5430 2090 5460
rect 2020 5390 2090 5430
rect 2020 5330 2040 5390
rect 2070 5330 2090 5390
rect 2020 5290 2090 5330
rect 2020 5230 2040 5290
rect 2070 5230 2090 5290
rect 2020 5190 2090 5230
rect 2020 5130 2040 5190
rect 2070 5130 2090 5190
rect 2020 5090 2090 5130
rect 2020 5030 2040 5090
rect 2070 5030 2090 5090
rect 2020 4990 2090 5030
rect 2020 4930 2040 4990
rect 2070 4930 2090 4990
rect 2020 4890 2090 4930
rect 2020 4830 2040 4890
rect 2070 4830 2090 4890
rect 2020 4790 2090 4830
rect 2020 4730 2040 4790
rect 2070 4730 2090 4790
rect 2020 4690 2090 4730
rect 2020 4630 2040 4690
rect 2070 4630 2090 4690
rect 2020 4590 2090 4630
rect 2020 4530 2040 4590
rect 2070 4530 2090 4590
rect 2020 4490 2090 4530
rect 2020 4460 2040 4490
rect 2070 4460 2090 4490
rect 2190 5430 2210 5460
rect 2240 5430 2260 5460
rect 2190 5390 2260 5430
rect 2190 5330 2210 5390
rect 2240 5330 2260 5390
rect 2190 5290 2260 5330
rect 2190 5230 2210 5290
rect 2240 5230 2260 5290
rect 2190 5190 2260 5230
rect 2190 5130 2210 5190
rect 2240 5130 2260 5190
rect 2190 5090 2260 5130
rect 2190 5030 2210 5090
rect 2240 5030 2260 5090
rect 2190 4990 2260 5030
rect 2190 4930 2210 4990
rect 2240 4930 2260 4990
rect 2190 4890 2260 4930
rect 2190 4830 2210 4890
rect 2240 4830 2260 4890
rect 2190 4790 2260 4830
rect 2190 4730 2210 4790
rect 2240 4730 2260 4790
rect 2190 4690 2260 4730
rect 2190 4630 2210 4690
rect 2240 4630 2260 4690
rect 2190 4590 2260 4630
rect 2190 4530 2210 4590
rect 2240 4530 2260 4590
rect 2190 4490 2260 4530
rect 2190 4460 2210 4490
rect 2240 4460 2260 4490
rect 2360 5430 2380 5460
rect 2410 5430 2430 5460
rect 2360 5390 2430 5430
rect 2360 5330 2380 5390
rect 2410 5330 2430 5390
rect 2360 5290 2430 5330
rect 2360 5230 2380 5290
rect 2410 5230 2430 5290
rect 2360 5190 2430 5230
rect 2360 5130 2380 5190
rect 2410 5130 2430 5190
rect 2360 5090 2430 5130
rect 2360 5030 2380 5090
rect 2410 5030 2430 5090
rect 2360 4990 2430 5030
rect 2360 4930 2380 4990
rect 2410 4930 2430 4990
rect 2360 4890 2430 4930
rect 2360 4830 2380 4890
rect 2410 4830 2430 4890
rect 2360 4790 2430 4830
rect 2360 4730 2380 4790
rect 2410 4730 2430 4790
rect 2360 4690 2430 4730
rect 2360 4630 2380 4690
rect 2410 4630 2430 4690
rect 2360 4590 2430 4630
rect 2360 4530 2380 4590
rect 2410 4530 2430 4590
rect 2360 4490 2430 4530
rect 2360 4460 2380 4490
rect 2410 4460 2430 4490
rect 2530 5430 2550 5460
rect 2580 5430 2600 5460
rect 2530 5390 2600 5430
rect 2530 5330 2550 5390
rect 2580 5330 2600 5390
rect 2530 5290 2600 5330
rect 2530 5230 2550 5290
rect 2580 5230 2600 5290
rect 2530 5190 2600 5230
rect 2530 5130 2550 5190
rect 2580 5130 2600 5190
rect 2530 5090 2600 5130
rect 2530 5030 2550 5090
rect 2580 5030 2600 5090
rect 2530 4990 2600 5030
rect 2530 4930 2550 4990
rect 2580 4930 2600 4990
rect 2530 4890 2600 4930
rect 2530 4830 2550 4890
rect 2580 4830 2600 4890
rect 2530 4790 2600 4830
rect 2530 4730 2550 4790
rect 2580 4730 2600 4790
rect 2530 4690 2600 4730
rect 2530 4630 2550 4690
rect 2580 4630 2600 4690
rect 2530 4590 2600 4630
rect 2530 4530 2550 4590
rect 2580 4530 2600 4590
rect 2530 4490 2600 4530
rect 2530 4460 2550 4490
rect 2580 4460 2600 4490
rect 2700 5430 2720 5460
rect 2750 5430 2770 5460
rect 2700 5390 2770 5430
rect 2700 5330 2720 5390
rect 2750 5330 2770 5390
rect 2700 5290 2770 5330
rect 2700 5230 2720 5290
rect 2750 5230 2770 5290
rect 2700 5190 2770 5230
rect 2700 5130 2720 5190
rect 2750 5130 2770 5190
rect 2700 5090 2770 5130
rect 2700 5030 2720 5090
rect 2750 5030 2770 5090
rect 2700 4990 2770 5030
rect 2700 4930 2720 4990
rect 2750 4930 2770 4990
rect 2700 4890 2770 4930
rect 2700 4830 2720 4890
rect 2750 4830 2770 4890
rect 2700 4790 2770 4830
rect 2700 4730 2720 4790
rect 2750 4730 2770 4790
rect 2700 4690 2770 4730
rect 2700 4630 2720 4690
rect 2750 4630 2770 4690
rect 2700 4590 2770 4630
rect 2700 4530 2720 4590
rect 2750 4530 2770 4590
rect 2700 4490 2770 4530
rect 2700 4460 2720 4490
rect 2750 4460 2770 4490
rect 2870 5430 2890 5460
rect 2920 5430 2940 5460
rect 2870 5390 2940 5430
rect 2870 5330 2890 5390
rect 2920 5330 2940 5390
rect 2870 5290 2940 5330
rect 2870 5230 2890 5290
rect 2920 5230 2940 5290
rect 2870 5190 2940 5230
rect 2870 5130 2890 5190
rect 2920 5130 2940 5190
rect 2870 5090 2940 5130
rect 2870 5030 2890 5090
rect 2920 5030 2940 5090
rect 2870 4990 2940 5030
rect 2870 4930 2890 4990
rect 2920 4930 2940 4990
rect 2870 4890 2940 4930
rect 2870 4830 2890 4890
rect 2920 4830 2940 4890
rect 2870 4790 2940 4830
rect 2870 4730 2890 4790
rect 2920 4730 2940 4790
rect 2870 4690 2940 4730
rect 2870 4630 2890 4690
rect 2920 4630 2940 4690
rect 2870 4590 2940 4630
rect 2870 4530 2890 4590
rect 2920 4530 2940 4590
rect 2870 4490 2940 4530
rect 2870 4460 2890 4490
rect 2920 4460 2940 4490
rect 3040 5430 3060 5460
rect 3090 5430 3110 5460
rect 3040 5390 3110 5430
rect 3040 5330 3060 5390
rect 3090 5330 3110 5390
rect 3040 5290 3110 5330
rect 3040 5230 3060 5290
rect 3090 5230 3110 5290
rect 3040 5190 3110 5230
rect 3040 5130 3060 5190
rect 3090 5130 3110 5190
rect 3040 5090 3110 5130
rect 3040 5030 3060 5090
rect 3090 5030 3110 5090
rect 3040 4990 3110 5030
rect 3040 4930 3060 4990
rect 3090 4930 3110 4990
rect 3040 4890 3110 4930
rect 3040 4830 3060 4890
rect 3090 4830 3110 4890
rect 3040 4790 3110 4830
rect 3040 4730 3060 4790
rect 3090 4730 3110 4790
rect 3040 4690 3110 4730
rect 3040 4630 3060 4690
rect 3090 4630 3110 4690
rect 3040 4590 3110 4630
rect 3040 4530 3060 4590
rect 3090 4530 3110 4590
rect 3040 4490 3110 4530
rect 3040 4460 3060 4490
rect 3090 4460 3110 4490
rect 3210 5430 3230 5460
rect 3260 5430 3280 5460
rect 3210 5390 3280 5430
rect 3210 5330 3230 5390
rect 3260 5330 3280 5390
rect 3210 5290 3280 5330
rect 3210 5230 3230 5290
rect 3260 5230 3280 5290
rect 3210 5190 3280 5230
rect 3210 5130 3230 5190
rect 3260 5130 3280 5190
rect 3210 5090 3280 5130
rect 3210 5030 3230 5090
rect 3260 5030 3280 5090
rect 3210 4990 3280 5030
rect 3210 4930 3230 4990
rect 3260 4930 3280 4990
rect 3210 4890 3280 4930
rect 3210 4830 3230 4890
rect 3260 4830 3280 4890
rect 3210 4790 3280 4830
rect 3210 4730 3230 4790
rect 3260 4730 3280 4790
rect 3210 4690 3280 4730
rect 3210 4630 3230 4690
rect 3260 4630 3280 4690
rect 3210 4590 3280 4630
rect 3210 4530 3230 4590
rect 3260 4530 3280 4590
rect 3210 4490 3280 4530
rect 3210 4460 3230 4490
rect 3260 4460 3280 4490
rect 3380 4460 3400 5460
rect 3440 5100 3460 5600
rect 3660 5100 3690 5600
rect 3430 4560 3460 5060
rect 3660 4560 3680 5060
rect 3430 4500 3450 4560
rect 3430 4490 3470 4500
rect 3430 4470 3440 4490
rect 3460 4470 3470 4490
rect 3430 4460 3470 4470
rect -210 4390 -60 4400
rect -210 4370 -200 4390
rect -180 4370 -60 4390
rect -210 4360 -60 4370
rect -160 4340 -60 4360
rect -20 4390 220 4400
rect -20 4370 90 4390
rect 110 4370 220 4390
rect -20 4360 220 4370
rect -20 4340 80 4360
rect 120 4340 220 4360
rect 260 4390 500 4400
rect 260 4370 370 4390
rect 390 4370 500 4390
rect 260 4360 500 4370
rect 260 4340 360 4360
rect 400 4340 500 4360
rect 540 4390 780 4400
rect 540 4370 650 4390
rect 670 4370 780 4390
rect 540 4360 780 4370
rect 540 4340 640 4360
rect 680 4340 780 4360
rect 820 4390 1060 4400
rect 820 4370 930 4390
rect 950 4370 1060 4390
rect 820 4360 1060 4370
rect 820 4340 920 4360
rect 960 4340 1060 4360
rect 1100 4390 1340 4400
rect 1100 4370 1210 4390
rect 1230 4370 1340 4390
rect 1100 4360 1340 4370
rect 1610 4390 1770 4400
rect 1610 4370 1620 4390
rect 1640 4370 1740 4390
rect 1760 4370 1770 4390
rect 1610 4360 1770 4370
rect 2040 4390 2280 4400
rect 2040 4370 2150 4390
rect 2170 4370 2280 4390
rect 2040 4360 2280 4370
rect 1100 4340 1200 4360
rect 1240 4340 1340 4360
rect 2040 4340 2140 4360
rect 2180 4340 2280 4360
rect 2320 4390 2560 4400
rect 2320 4370 2430 4390
rect 2450 4370 2560 4390
rect 2320 4360 2560 4370
rect 2320 4340 2420 4360
rect 2460 4340 2560 4360
rect 2600 4390 2840 4400
rect 2600 4370 2710 4390
rect 2730 4370 2840 4390
rect 2600 4360 2840 4370
rect 2600 4340 2700 4360
rect 2740 4340 2840 4360
rect 2880 4390 3120 4400
rect 2880 4370 2990 4390
rect 3010 4370 3120 4390
rect 2880 4360 3120 4370
rect 2880 4340 2980 4360
rect 3020 4340 3120 4360
rect 3160 4390 3400 4400
rect 3160 4370 3270 4390
rect 3290 4370 3400 4390
rect 3160 4360 3400 4370
rect 3160 4340 3260 4360
rect 3300 4340 3400 4360
rect 3440 4390 3590 4400
rect 3440 4370 3560 4390
rect 3580 4370 3590 4390
rect 3440 4360 3590 4370
rect 3440 4340 3540 4360
rect -160 3300 -60 3340
rect -20 3300 80 3340
rect 120 3300 220 3340
rect 260 3300 360 3340
rect 400 3300 500 3340
rect 540 3300 640 3340
rect 680 3300 780 3340
rect 820 3300 920 3340
rect 960 3300 1060 3340
rect 1100 3300 1200 3340
rect 1240 3300 1340 3340
rect 2040 3300 2140 3340
rect 2180 3300 2280 3340
rect 2320 3300 2420 3340
rect 2460 3300 2560 3340
rect 2600 3300 2700 3340
rect 2740 3300 2840 3340
rect 2880 3300 2980 3340
rect 3020 3300 3120 3340
rect 3160 3300 3260 3340
rect 3300 3300 3400 3340
rect 3440 3300 3540 3340
rect -160 2280 -60 2300
rect -210 2270 -60 2280
rect -210 2250 -200 2270
rect -180 2250 -60 2270
rect -210 2240 -60 2250
rect -20 2280 80 2300
rect 120 2280 220 2300
rect -20 2270 220 2280
rect -20 2250 90 2270
rect 110 2250 220 2270
rect -20 2240 220 2250
rect 260 2280 360 2300
rect 400 2280 500 2300
rect 260 2270 500 2280
rect 260 2250 370 2270
rect 390 2250 500 2270
rect 260 2240 500 2250
rect 540 2280 640 2300
rect 680 2280 780 2300
rect 540 2270 780 2280
rect 540 2250 650 2270
rect 670 2250 780 2270
rect 540 2240 780 2250
rect 820 2280 920 2300
rect 960 2280 1060 2300
rect 820 2270 1060 2280
rect 820 2250 930 2270
rect 950 2250 1060 2270
rect 820 2240 1060 2250
rect 1100 2280 1200 2300
rect 1240 2280 1340 2300
rect 2040 2280 2140 2300
rect 2180 2280 2280 2300
rect 1100 2270 1340 2280
rect 1100 2250 1210 2270
rect 1230 2250 1340 2270
rect 1100 2240 1340 2250
rect 1610 2270 1770 2280
rect 1610 2250 1620 2270
rect 1640 2250 1740 2270
rect 1760 2250 1770 2270
rect 1610 2240 1770 2250
rect 2040 2270 2280 2280
rect 2040 2250 2150 2270
rect 2170 2250 2280 2270
rect 2040 2240 2280 2250
rect 2320 2280 2420 2300
rect 2460 2280 2560 2300
rect 2320 2270 2560 2280
rect 2320 2250 2430 2270
rect 2450 2250 2560 2270
rect 2320 2240 2560 2250
rect 2600 2280 2700 2300
rect 2740 2280 2840 2300
rect 2600 2270 2840 2280
rect 2600 2250 2710 2270
rect 2730 2250 2840 2270
rect 2600 2240 2840 2250
rect 2880 2280 2980 2300
rect 3020 2280 3120 2300
rect 2880 2270 3120 2280
rect 2880 2250 2990 2270
rect 3010 2250 3120 2270
rect 2880 2240 3120 2250
rect 3160 2280 3260 2300
rect 3300 2280 3400 2300
rect 3160 2270 3400 2280
rect 3160 2250 3270 2270
rect 3290 2250 3400 2270
rect 3160 2240 3400 2250
rect 3440 2280 3540 2300
rect 3440 2270 3590 2280
rect 3440 2250 3560 2270
rect 3580 2250 3590 2270
rect 3440 2240 3590 2250
rect -90 2170 -50 2180
rect -90 2150 -80 2170
rect -60 2150 -50 2170
rect -90 2140 -50 2150
rect -70 2080 -50 2140
rect -300 1580 -280 2080
rect -80 1580 -50 2080
rect -310 1040 -280 1540
rect -80 1040 -60 1540
rect -20 1180 0 2180
rect 100 2150 120 2180
rect 150 2150 170 2180
rect 100 2110 170 2150
rect 100 2050 120 2110
rect 150 2050 170 2110
rect 100 2010 170 2050
rect 100 1950 120 2010
rect 150 1950 170 2010
rect 100 1910 170 1950
rect 100 1850 120 1910
rect 150 1850 170 1910
rect 100 1810 170 1850
rect 100 1750 120 1810
rect 150 1750 170 1810
rect 100 1710 170 1750
rect 100 1650 120 1710
rect 150 1650 170 1710
rect 100 1610 170 1650
rect 100 1550 120 1610
rect 150 1550 170 1610
rect 100 1510 170 1550
rect 100 1450 120 1510
rect 150 1450 170 1510
rect 100 1410 170 1450
rect 100 1350 120 1410
rect 150 1350 170 1410
rect 100 1310 170 1350
rect 100 1250 120 1310
rect 150 1250 170 1310
rect 100 1210 170 1250
rect 100 1180 120 1210
rect 150 1180 170 1210
rect 270 2150 290 2180
rect 320 2150 340 2180
rect 270 2110 340 2150
rect 270 2050 290 2110
rect 320 2050 340 2110
rect 270 2010 340 2050
rect 270 1950 290 2010
rect 320 1950 340 2010
rect 270 1910 340 1950
rect 270 1850 290 1910
rect 320 1850 340 1910
rect 270 1810 340 1850
rect 270 1750 290 1810
rect 320 1750 340 1810
rect 270 1710 340 1750
rect 270 1650 290 1710
rect 320 1650 340 1710
rect 270 1610 340 1650
rect 270 1550 290 1610
rect 320 1550 340 1610
rect 270 1510 340 1550
rect 270 1450 290 1510
rect 320 1450 340 1510
rect 270 1410 340 1450
rect 270 1350 290 1410
rect 320 1350 340 1410
rect 270 1310 340 1350
rect 270 1250 290 1310
rect 320 1250 340 1310
rect 270 1210 340 1250
rect 270 1180 290 1210
rect 320 1180 340 1210
rect 440 2150 460 2180
rect 490 2150 510 2180
rect 440 2110 510 2150
rect 440 2050 460 2110
rect 490 2050 510 2110
rect 440 2010 510 2050
rect 440 1950 460 2010
rect 490 1950 510 2010
rect 440 1910 510 1950
rect 440 1850 460 1910
rect 490 1850 510 1910
rect 440 1810 510 1850
rect 440 1750 460 1810
rect 490 1750 510 1810
rect 440 1710 510 1750
rect 440 1650 460 1710
rect 490 1650 510 1710
rect 440 1610 510 1650
rect 440 1550 460 1610
rect 490 1550 510 1610
rect 440 1510 510 1550
rect 440 1450 460 1510
rect 490 1450 510 1510
rect 440 1410 510 1450
rect 440 1350 460 1410
rect 490 1350 510 1410
rect 440 1310 510 1350
rect 440 1250 460 1310
rect 490 1250 510 1310
rect 440 1210 510 1250
rect 440 1180 460 1210
rect 490 1180 510 1210
rect 610 2150 630 2180
rect 660 2150 680 2180
rect 610 2110 680 2150
rect 610 2050 630 2110
rect 660 2050 680 2110
rect 610 2010 680 2050
rect 610 1950 630 2010
rect 660 1950 680 2010
rect 610 1910 680 1950
rect 610 1850 630 1910
rect 660 1850 680 1910
rect 610 1810 680 1850
rect 610 1750 630 1810
rect 660 1750 680 1810
rect 610 1710 680 1750
rect 610 1650 630 1710
rect 660 1650 680 1710
rect 610 1610 680 1650
rect 610 1550 630 1610
rect 660 1550 680 1610
rect 610 1510 680 1550
rect 610 1450 630 1510
rect 660 1450 680 1510
rect 610 1410 680 1450
rect 610 1350 630 1410
rect 660 1350 680 1410
rect 610 1310 680 1350
rect 610 1250 630 1310
rect 660 1250 680 1310
rect 610 1210 680 1250
rect 610 1180 630 1210
rect 660 1180 680 1210
rect 780 2150 800 2180
rect 830 2150 850 2180
rect 780 2110 850 2150
rect 780 2050 800 2110
rect 830 2050 850 2110
rect 780 2010 850 2050
rect 780 1950 800 2010
rect 830 1950 850 2010
rect 780 1910 850 1950
rect 780 1850 800 1910
rect 830 1850 850 1910
rect 780 1810 850 1850
rect 780 1750 800 1810
rect 830 1750 850 1810
rect 780 1710 850 1750
rect 780 1650 800 1710
rect 830 1650 850 1710
rect 780 1610 850 1650
rect 780 1550 800 1610
rect 830 1550 850 1610
rect 780 1510 850 1550
rect 780 1450 800 1510
rect 830 1450 850 1510
rect 780 1410 850 1450
rect 780 1350 800 1410
rect 830 1350 850 1410
rect 780 1310 850 1350
rect 780 1250 800 1310
rect 830 1250 850 1310
rect 780 1210 850 1250
rect 780 1180 800 1210
rect 830 1180 850 1210
rect 950 2150 970 2180
rect 1000 2150 1020 2180
rect 950 2110 1020 2150
rect 950 2050 970 2110
rect 1000 2050 1020 2110
rect 950 2010 1020 2050
rect 950 1950 970 2010
rect 1000 1950 1020 2010
rect 950 1910 1020 1950
rect 950 1850 970 1910
rect 1000 1850 1020 1910
rect 950 1810 1020 1850
rect 950 1750 970 1810
rect 1000 1750 1020 1810
rect 950 1710 1020 1750
rect 950 1650 970 1710
rect 1000 1650 1020 1710
rect 950 1610 1020 1650
rect 950 1550 970 1610
rect 1000 1550 1020 1610
rect 950 1510 1020 1550
rect 950 1450 970 1510
rect 1000 1450 1020 1510
rect 950 1410 1020 1450
rect 950 1350 970 1410
rect 1000 1350 1020 1410
rect 950 1310 1020 1350
rect 950 1250 970 1310
rect 1000 1250 1020 1310
rect 950 1210 1020 1250
rect 950 1180 970 1210
rect 1000 1180 1020 1210
rect 1120 2150 1140 2180
rect 1170 2150 1190 2180
rect 1120 2110 1190 2150
rect 1120 2050 1140 2110
rect 1170 2050 1190 2110
rect 1120 2010 1190 2050
rect 1120 1950 1140 2010
rect 1170 1950 1190 2010
rect 1120 1910 1190 1950
rect 1120 1850 1140 1910
rect 1170 1850 1190 1910
rect 1120 1810 1190 1850
rect 1120 1750 1140 1810
rect 1170 1750 1190 1810
rect 1120 1710 1190 1750
rect 1120 1650 1140 1710
rect 1170 1650 1190 1710
rect 1120 1610 1190 1650
rect 1120 1550 1140 1610
rect 1170 1550 1190 1610
rect 1120 1510 1190 1550
rect 1120 1450 1140 1510
rect 1170 1450 1190 1510
rect 1120 1410 1190 1450
rect 1120 1350 1140 1410
rect 1170 1350 1190 1410
rect 1120 1310 1190 1350
rect 1120 1250 1140 1310
rect 1170 1250 1190 1310
rect 1120 1210 1190 1250
rect 1120 1180 1140 1210
rect 1170 1180 1190 1210
rect 1290 2150 1310 2180
rect 1340 2150 1360 2180
rect 1290 2110 1360 2150
rect 1290 2050 1310 2110
rect 1340 2050 1360 2110
rect 1290 2010 1360 2050
rect 1290 1950 1310 2010
rect 1340 1950 1360 2010
rect 1290 1910 1360 1950
rect 1290 1850 1310 1910
rect 1340 1850 1360 1910
rect 1290 1810 1360 1850
rect 1290 1750 1310 1810
rect 1340 1750 1360 1810
rect 1290 1710 1360 1750
rect 1290 1650 1310 1710
rect 1340 1650 1360 1710
rect 1290 1610 1360 1650
rect 1290 1550 1310 1610
rect 1340 1550 1360 1610
rect 1290 1510 1360 1550
rect 1290 1450 1310 1510
rect 1340 1450 1360 1510
rect 1290 1410 1360 1450
rect 1290 1350 1310 1410
rect 1340 1350 1360 1410
rect 1290 1310 1360 1350
rect 1290 1250 1310 1310
rect 1340 1250 1360 1310
rect 1290 1210 1360 1250
rect 1290 1180 1310 1210
rect 1340 1180 1360 1210
rect 1460 2150 1480 2180
rect 1510 2150 1530 2180
rect 1460 2110 1530 2150
rect 1460 2050 1480 2110
rect 1510 2050 1530 2110
rect 1460 2010 1530 2050
rect 1460 1950 1480 2010
rect 1510 1950 1530 2010
rect 1460 1910 1530 1950
rect 1460 1850 1480 1910
rect 1510 1850 1530 1910
rect 1460 1810 1530 1850
rect 1460 1750 1480 1810
rect 1510 1750 1530 1810
rect 1460 1710 1530 1750
rect 1460 1650 1480 1710
rect 1510 1650 1530 1710
rect 1460 1610 1530 1650
rect 1460 1550 1480 1610
rect 1510 1550 1530 1610
rect 1460 1510 1530 1550
rect 1460 1450 1480 1510
rect 1510 1450 1530 1510
rect 1460 1410 1530 1450
rect 1460 1350 1480 1410
rect 1510 1350 1530 1410
rect 1460 1310 1530 1350
rect 1460 1250 1480 1310
rect 1510 1250 1530 1310
rect 1460 1210 1530 1250
rect 1460 1180 1480 1210
rect 1510 1180 1530 1210
rect 1630 2150 1650 2180
rect 1680 2150 1700 2240
rect 1730 2150 1750 2180
rect 1630 2110 1750 2150
rect 1630 2050 1650 2110
rect 1680 2050 1700 2110
rect 1730 2050 1750 2110
rect 1630 2010 1750 2050
rect 1630 1950 1650 2010
rect 1680 1950 1700 2010
rect 1730 1950 1750 2010
rect 1630 1910 1750 1950
rect 1630 1850 1650 1910
rect 1680 1850 1700 1910
rect 1730 1850 1750 1910
rect 1630 1810 1750 1850
rect 1630 1750 1650 1810
rect 1680 1750 1700 1810
rect 1730 1750 1750 1810
rect 1630 1710 1750 1750
rect 1630 1650 1650 1710
rect 1680 1650 1700 1710
rect 1730 1650 1750 1710
rect 1630 1610 1750 1650
rect 1630 1550 1650 1610
rect 1680 1550 1700 1610
rect 1730 1550 1750 1610
rect 1630 1510 1750 1550
rect 1630 1450 1650 1510
rect 1680 1450 1700 1510
rect 1730 1450 1750 1510
rect 1630 1410 1750 1450
rect 1630 1350 1650 1410
rect 1680 1350 1700 1410
rect 1730 1350 1750 1410
rect 1630 1310 1750 1350
rect 1630 1250 1650 1310
rect 1680 1250 1700 1310
rect 1730 1250 1750 1310
rect 1630 1210 1750 1250
rect 1630 1180 1650 1210
rect -20 1040 0 1140
rect 100 1110 120 1140
rect 150 1110 170 1140
rect 100 1070 170 1110
rect 100 1040 120 1070
rect 150 1040 170 1070
rect 270 1110 290 1140
rect 320 1110 340 1140
rect 270 1070 340 1110
rect 270 1040 290 1070
rect 320 1040 340 1070
rect 440 1110 460 1140
rect 490 1110 510 1140
rect 440 1070 510 1110
rect 440 1040 460 1070
rect 490 1040 510 1070
rect 610 1110 630 1140
rect 660 1110 680 1140
rect 610 1070 680 1110
rect 610 1040 630 1070
rect 660 1040 680 1070
rect 780 1110 800 1140
rect 830 1110 850 1140
rect 780 1070 850 1110
rect 780 1040 800 1070
rect 830 1040 850 1070
rect 950 1110 970 1140
rect 1000 1110 1020 1140
rect 950 1070 1020 1110
rect 950 1040 970 1070
rect 1000 1040 1020 1070
rect 1120 1110 1140 1140
rect 1170 1110 1190 1140
rect 1120 1070 1190 1110
rect 1120 1040 1140 1070
rect 1170 1040 1190 1070
rect 1290 1110 1310 1140
rect 1340 1110 1360 1140
rect 1290 1070 1360 1110
rect 1290 1040 1310 1070
rect 1340 1040 1360 1070
rect 1460 1110 1480 1140
rect 1510 1110 1530 1140
rect 1460 1070 1530 1110
rect 1460 1040 1480 1070
rect 1510 1040 1530 1070
rect 1630 1110 1650 1140
rect 1680 1110 1700 1210
rect 1730 1180 1750 1210
rect 1850 2150 1870 2180
rect 1900 2150 1920 2180
rect 1850 2110 1920 2150
rect 1850 2050 1870 2110
rect 1900 2050 1920 2110
rect 1850 2010 1920 2050
rect 1850 1950 1870 2010
rect 1900 1950 1920 2010
rect 1850 1910 1920 1950
rect 1850 1850 1870 1910
rect 1900 1850 1920 1910
rect 1850 1810 1920 1850
rect 1850 1750 1870 1810
rect 1900 1750 1920 1810
rect 1850 1710 1920 1750
rect 1850 1650 1870 1710
rect 1900 1650 1920 1710
rect 1850 1610 1920 1650
rect 1850 1550 1870 1610
rect 1900 1550 1920 1610
rect 1850 1510 1920 1550
rect 1850 1450 1870 1510
rect 1900 1450 1920 1510
rect 1850 1410 1920 1450
rect 1850 1350 1870 1410
rect 1900 1350 1920 1410
rect 1850 1310 1920 1350
rect 1850 1250 1870 1310
rect 1900 1250 1920 1310
rect 1850 1210 1920 1250
rect 1850 1180 1870 1210
rect 1900 1180 1920 1210
rect 2020 2150 2040 2180
rect 2070 2150 2090 2180
rect 2020 2110 2090 2150
rect 2020 2050 2040 2110
rect 2070 2050 2090 2110
rect 2020 2010 2090 2050
rect 2020 1950 2040 2010
rect 2070 1950 2090 2010
rect 2020 1910 2090 1950
rect 2020 1850 2040 1910
rect 2070 1850 2090 1910
rect 2020 1810 2090 1850
rect 2020 1750 2040 1810
rect 2070 1750 2090 1810
rect 2020 1710 2090 1750
rect 2020 1650 2040 1710
rect 2070 1650 2090 1710
rect 2020 1610 2090 1650
rect 2020 1550 2040 1610
rect 2070 1550 2090 1610
rect 2020 1510 2090 1550
rect 2020 1450 2040 1510
rect 2070 1450 2090 1510
rect 2020 1410 2090 1450
rect 2020 1350 2040 1410
rect 2070 1350 2090 1410
rect 2020 1310 2090 1350
rect 2020 1250 2040 1310
rect 2070 1250 2090 1310
rect 2020 1210 2090 1250
rect 2020 1180 2040 1210
rect 2070 1180 2090 1210
rect 2190 2150 2210 2180
rect 2240 2150 2260 2180
rect 2190 2110 2260 2150
rect 2190 2050 2210 2110
rect 2240 2050 2260 2110
rect 2190 2010 2260 2050
rect 2190 1950 2210 2010
rect 2240 1950 2260 2010
rect 2190 1910 2260 1950
rect 2190 1850 2210 1910
rect 2240 1850 2260 1910
rect 2190 1810 2260 1850
rect 2190 1750 2210 1810
rect 2240 1750 2260 1810
rect 2190 1710 2260 1750
rect 2190 1650 2210 1710
rect 2240 1650 2260 1710
rect 2190 1610 2260 1650
rect 2190 1550 2210 1610
rect 2240 1550 2260 1610
rect 2190 1510 2260 1550
rect 2190 1450 2210 1510
rect 2240 1450 2260 1510
rect 2190 1410 2260 1450
rect 2190 1350 2210 1410
rect 2240 1350 2260 1410
rect 2190 1310 2260 1350
rect 2190 1250 2210 1310
rect 2240 1250 2260 1310
rect 2190 1210 2260 1250
rect 2190 1180 2210 1210
rect 2240 1180 2260 1210
rect 2360 2150 2380 2180
rect 2410 2150 2430 2180
rect 2360 2110 2430 2150
rect 2360 2050 2380 2110
rect 2410 2050 2430 2110
rect 2360 2010 2430 2050
rect 2360 1950 2380 2010
rect 2410 1950 2430 2010
rect 2360 1910 2430 1950
rect 2360 1850 2380 1910
rect 2410 1850 2430 1910
rect 2360 1810 2430 1850
rect 2360 1750 2380 1810
rect 2410 1750 2430 1810
rect 2360 1710 2430 1750
rect 2360 1650 2380 1710
rect 2410 1650 2430 1710
rect 2360 1610 2430 1650
rect 2360 1550 2380 1610
rect 2410 1550 2430 1610
rect 2360 1510 2430 1550
rect 2360 1450 2380 1510
rect 2410 1450 2430 1510
rect 2360 1410 2430 1450
rect 2360 1350 2380 1410
rect 2410 1350 2430 1410
rect 2360 1310 2430 1350
rect 2360 1250 2380 1310
rect 2410 1250 2430 1310
rect 2360 1210 2430 1250
rect 2360 1180 2380 1210
rect 2410 1180 2430 1210
rect 2530 2150 2550 2180
rect 2580 2150 2600 2180
rect 2530 2110 2600 2150
rect 2530 2050 2550 2110
rect 2580 2050 2600 2110
rect 2530 2010 2600 2050
rect 2530 1950 2550 2010
rect 2580 1950 2600 2010
rect 2530 1910 2600 1950
rect 2530 1850 2550 1910
rect 2580 1850 2600 1910
rect 2530 1810 2600 1850
rect 2530 1750 2550 1810
rect 2580 1750 2600 1810
rect 2530 1710 2600 1750
rect 2530 1650 2550 1710
rect 2580 1650 2600 1710
rect 2530 1610 2600 1650
rect 2530 1550 2550 1610
rect 2580 1550 2600 1610
rect 2530 1510 2600 1550
rect 2530 1450 2550 1510
rect 2580 1450 2600 1510
rect 2530 1410 2600 1450
rect 2530 1350 2550 1410
rect 2580 1350 2600 1410
rect 2530 1310 2600 1350
rect 2530 1250 2550 1310
rect 2580 1250 2600 1310
rect 2530 1210 2600 1250
rect 2530 1180 2550 1210
rect 2580 1180 2600 1210
rect 2700 2150 2720 2180
rect 2750 2150 2770 2180
rect 2700 2110 2770 2150
rect 2700 2050 2720 2110
rect 2750 2050 2770 2110
rect 2700 2010 2770 2050
rect 2700 1950 2720 2010
rect 2750 1950 2770 2010
rect 2700 1910 2770 1950
rect 2700 1850 2720 1910
rect 2750 1850 2770 1910
rect 2700 1810 2770 1850
rect 2700 1750 2720 1810
rect 2750 1750 2770 1810
rect 2700 1710 2770 1750
rect 2700 1650 2720 1710
rect 2750 1650 2770 1710
rect 2700 1610 2770 1650
rect 2700 1550 2720 1610
rect 2750 1550 2770 1610
rect 2700 1510 2770 1550
rect 2700 1450 2720 1510
rect 2750 1450 2770 1510
rect 2700 1410 2770 1450
rect 2700 1350 2720 1410
rect 2750 1350 2770 1410
rect 2700 1310 2770 1350
rect 2700 1250 2720 1310
rect 2750 1250 2770 1310
rect 2700 1210 2770 1250
rect 2700 1180 2720 1210
rect 2750 1180 2770 1210
rect 2870 2150 2890 2180
rect 2920 2150 2940 2180
rect 2870 2110 2940 2150
rect 2870 2050 2890 2110
rect 2920 2050 2940 2110
rect 2870 2010 2940 2050
rect 2870 1950 2890 2010
rect 2920 1950 2940 2010
rect 2870 1910 2940 1950
rect 2870 1850 2890 1910
rect 2920 1850 2940 1910
rect 2870 1810 2940 1850
rect 2870 1750 2890 1810
rect 2920 1750 2940 1810
rect 2870 1710 2940 1750
rect 2870 1650 2890 1710
rect 2920 1650 2940 1710
rect 2870 1610 2940 1650
rect 2870 1550 2890 1610
rect 2920 1550 2940 1610
rect 2870 1510 2940 1550
rect 2870 1450 2890 1510
rect 2920 1450 2940 1510
rect 2870 1410 2940 1450
rect 2870 1350 2890 1410
rect 2920 1350 2940 1410
rect 2870 1310 2940 1350
rect 2870 1250 2890 1310
rect 2920 1250 2940 1310
rect 2870 1210 2940 1250
rect 2870 1180 2890 1210
rect 2920 1180 2940 1210
rect 3040 2150 3060 2180
rect 3090 2150 3110 2180
rect 3040 2110 3110 2150
rect 3040 2050 3060 2110
rect 3090 2050 3110 2110
rect 3040 2010 3110 2050
rect 3040 1950 3060 2010
rect 3090 1950 3110 2010
rect 3040 1910 3110 1950
rect 3040 1850 3060 1910
rect 3090 1850 3110 1910
rect 3040 1810 3110 1850
rect 3040 1750 3060 1810
rect 3090 1750 3110 1810
rect 3040 1710 3110 1750
rect 3040 1650 3060 1710
rect 3090 1650 3110 1710
rect 3040 1610 3110 1650
rect 3040 1550 3060 1610
rect 3090 1550 3110 1610
rect 3040 1510 3110 1550
rect 3040 1450 3060 1510
rect 3090 1450 3110 1510
rect 3040 1410 3110 1450
rect 3040 1350 3060 1410
rect 3090 1350 3110 1410
rect 3040 1310 3110 1350
rect 3040 1250 3060 1310
rect 3090 1250 3110 1310
rect 3040 1210 3110 1250
rect 3040 1180 3060 1210
rect 3090 1180 3110 1210
rect 3210 2150 3230 2180
rect 3260 2150 3280 2180
rect 3210 2110 3280 2150
rect 3210 2050 3230 2110
rect 3260 2050 3280 2110
rect 3210 2010 3280 2050
rect 3210 1950 3230 2010
rect 3260 1950 3280 2010
rect 3210 1910 3280 1950
rect 3210 1850 3230 1910
rect 3260 1850 3280 1910
rect 3210 1810 3280 1850
rect 3210 1750 3230 1810
rect 3260 1750 3280 1810
rect 3210 1710 3280 1750
rect 3210 1650 3230 1710
rect 3260 1650 3280 1710
rect 3210 1610 3280 1650
rect 3210 1550 3230 1610
rect 3260 1550 3280 1610
rect 3210 1510 3280 1550
rect 3210 1450 3230 1510
rect 3260 1450 3280 1510
rect 3210 1410 3280 1450
rect 3210 1350 3230 1410
rect 3260 1350 3280 1410
rect 3210 1310 3280 1350
rect 3210 1250 3230 1310
rect 3260 1250 3280 1310
rect 3210 1210 3280 1250
rect 3210 1180 3230 1210
rect 3260 1180 3280 1210
rect 3380 1180 3400 2180
rect 3430 2170 3470 2180
rect 3430 2150 3440 2170
rect 3460 2150 3470 2170
rect 3430 2140 3470 2150
rect 3430 2080 3450 2140
rect 3430 1580 3460 2080
rect 3660 1580 3680 2080
rect 1730 1110 1750 1140
rect 1630 1070 1750 1110
rect 1630 1040 1650 1070
rect 1730 1040 1750 1070
rect 1850 1110 1870 1140
rect 1900 1110 1920 1140
rect 1850 1070 1920 1110
rect 1850 1040 1870 1070
rect 1900 1040 1920 1070
rect 2020 1110 2040 1140
rect 2070 1110 2090 1140
rect 2020 1070 2090 1110
rect 2020 1040 2040 1070
rect 2070 1040 2090 1070
rect 2190 1110 2210 1140
rect 2240 1110 2260 1140
rect 2190 1070 2260 1110
rect 2190 1040 2210 1070
rect 2240 1040 2260 1070
rect 2360 1110 2380 1140
rect 2410 1110 2430 1140
rect 2360 1070 2430 1110
rect 2360 1040 2380 1070
rect 2410 1040 2430 1070
rect 2530 1110 2550 1140
rect 2580 1110 2600 1140
rect 2530 1070 2600 1110
rect 2530 1040 2550 1070
rect 2580 1040 2600 1070
rect 2700 1110 2720 1140
rect 2750 1110 2770 1140
rect 2700 1070 2770 1110
rect 2700 1040 2720 1070
rect 2750 1040 2770 1070
rect 2870 1110 2890 1140
rect 2920 1110 2940 1140
rect 2870 1070 2940 1110
rect 2870 1040 2890 1070
rect 2920 1040 2940 1070
rect 3040 1110 3060 1140
rect 3090 1110 3110 1140
rect 3040 1070 3110 1110
rect 3040 1040 3060 1070
rect 3090 1040 3110 1070
rect 3210 1110 3230 1140
rect 3260 1110 3280 1140
rect 3210 1070 3280 1110
rect 3210 1040 3230 1070
rect 3260 1040 3280 1070
rect 3380 1040 3400 1140
rect 3440 1040 3460 1540
rect 3660 1040 3690 1540
rect -310 980 -290 1040
rect -310 970 -270 980
rect -310 950 -300 970
rect -280 950 -270 970
rect -310 940 -270 950
rect -60 900 0 1000
rect 100 970 120 1000
rect 150 970 170 1000
rect 100 930 170 970
rect 100 900 120 930
rect 150 900 170 930
rect 270 970 290 1000
rect 320 970 340 1000
rect 270 930 340 970
rect 270 900 290 930
rect 320 900 340 930
rect 440 970 460 1000
rect 490 970 510 1000
rect 440 930 510 970
rect 440 900 460 930
rect 490 900 510 930
rect 610 970 630 1000
rect 660 970 680 1000
rect 610 930 680 970
rect 610 900 630 930
rect 660 900 680 930
rect 780 970 800 1000
rect 830 970 850 1000
rect 780 930 850 970
rect 780 900 800 930
rect 830 900 850 930
rect 950 970 970 1000
rect 1000 970 1020 1000
rect 950 930 1020 970
rect 950 900 970 930
rect 1000 900 1020 930
rect 1120 970 1140 1000
rect 1170 970 1190 1000
rect 1120 930 1190 970
rect 1120 900 1140 930
rect 1170 900 1190 930
rect 1290 970 1310 1000
rect 1340 970 1360 1000
rect 1290 930 1360 970
rect 1290 900 1310 930
rect 1340 900 1360 930
rect 1460 970 1480 1000
rect 1510 970 1530 1000
rect 1460 930 1530 970
rect 1460 900 1480 930
rect 1510 900 1530 930
rect 1630 970 1650 1000
rect 1730 970 1750 1000
rect 1630 930 1750 970
rect 1630 900 1650 930
rect 1730 900 1750 930
rect 1850 970 1870 1000
rect 1900 970 1920 1000
rect 1850 930 1920 970
rect 1850 900 1870 930
rect 1900 900 1920 930
rect 2020 970 2040 1000
rect 2070 970 2090 1000
rect 2020 930 2090 970
rect 2020 900 2040 930
rect 2070 900 2090 930
rect 2190 970 2210 1000
rect 2240 970 2260 1000
rect 2190 930 2260 970
rect 2190 900 2210 930
rect 2240 900 2260 930
rect 2360 970 2380 1000
rect 2410 970 2430 1000
rect 2360 930 2430 970
rect 2360 900 2380 930
rect 2410 900 2430 930
rect 2530 970 2550 1000
rect 2580 970 2600 1000
rect 2530 930 2600 970
rect 2530 900 2550 930
rect 2580 900 2600 930
rect 2700 970 2720 1000
rect 2750 970 2770 1000
rect 2700 930 2770 970
rect 2700 900 2720 930
rect 2750 900 2770 930
rect 2870 970 2890 1000
rect 2920 970 2940 1000
rect 2870 930 2940 970
rect 2870 900 2890 930
rect 2920 900 2940 930
rect 3040 970 3060 1000
rect 3090 970 3110 1000
rect 3040 930 3110 970
rect 3040 900 3060 930
rect 3090 900 3110 930
rect 3210 970 3230 1000
rect 3260 970 3280 1000
rect 3210 930 3280 970
rect 3210 900 3230 930
rect 3260 900 3280 930
rect 3380 900 3440 1000
rect 3670 980 3690 1040
rect 3650 970 3690 980
rect 3650 950 3660 970
rect 3680 950 3690 970
rect 3650 940 3690 950
rect -60 870 -20 900
rect -60 850 -50 870
rect -30 850 -20 870
rect -60 840 -20 850
rect 3400 870 3440 900
rect 3400 850 3410 870
rect 3430 850 3440 870
rect 3400 840 3440 850
<< polycont >>
rect -50 5770 -30 5790
rect 3410 5770 3430 5790
rect -300 5670 -280 5690
rect 3660 5670 3680 5690
rect -80 4470 -60 4490
rect 3440 4470 3460 4490
rect -200 4370 -180 4390
rect 90 4370 110 4390
rect 370 4370 390 4390
rect 650 4370 670 4390
rect 930 4370 950 4390
rect 1210 4370 1230 4390
rect 1620 4370 1640 4390
rect 1740 4370 1760 4390
rect 2150 4370 2170 4390
rect 2430 4370 2450 4390
rect 2710 4370 2730 4390
rect 2990 4370 3010 4390
rect 3270 4370 3290 4390
rect 3560 4370 3580 4390
rect -200 2250 -180 2270
rect 90 2250 110 2270
rect 370 2250 390 2270
rect 650 2250 670 2270
rect 930 2250 950 2270
rect 1210 2250 1230 2270
rect 1620 2250 1640 2270
rect 1740 2250 1760 2270
rect 2150 2250 2170 2270
rect 2430 2250 2450 2270
rect 2710 2250 2730 2270
rect 2990 2250 3010 2270
rect 3270 2250 3290 2270
rect 3560 2250 3580 2270
rect -80 2150 -60 2170
rect 3440 2150 3460 2170
rect -300 950 -280 970
rect 3660 950 3680 970
rect -50 850 -30 870
rect 3410 850 3430 870
<< locali >>
rect 20 5800 30 5810
rect -60 5790 30 5800
rect 70 5800 80 5810
rect 190 5800 200 5810
rect 70 5790 200 5800
rect 240 5800 250 5810
rect 360 5800 370 5810
rect 240 5790 370 5800
rect 410 5800 420 5810
rect 530 5800 540 5810
rect 410 5790 540 5800
rect 580 5800 590 5810
rect 700 5800 710 5810
rect 580 5790 710 5800
rect 750 5800 760 5810
rect 870 5800 880 5810
rect 750 5790 880 5800
rect 920 5800 930 5810
rect 1040 5800 1050 5810
rect 920 5790 1050 5800
rect 1090 5800 1100 5810
rect 1210 5800 1220 5810
rect 1090 5790 1220 5800
rect 1260 5800 1270 5810
rect 1380 5800 1390 5810
rect 1260 5790 1390 5800
rect 1430 5800 1440 5810
rect 1550 5800 1560 5810
rect 1430 5790 1560 5800
rect 1600 5800 1610 5810
rect 1770 5800 1780 5810
rect 1600 5790 1780 5800
rect 1820 5800 1830 5810
rect 1940 5800 1950 5810
rect 1820 5790 1950 5800
rect 1990 5800 2000 5810
rect 2110 5800 2120 5810
rect 1990 5790 2120 5800
rect 2160 5800 2170 5810
rect 2280 5800 2290 5810
rect 2160 5790 2290 5800
rect 2330 5800 2340 5810
rect 2450 5800 2460 5810
rect 2330 5790 2460 5800
rect 2500 5800 2510 5810
rect 2620 5800 2630 5810
rect 2500 5790 2630 5800
rect 2670 5800 2680 5810
rect 2790 5800 2800 5810
rect 2670 5790 2800 5800
rect 2840 5800 2850 5810
rect 2960 5800 2970 5810
rect 2840 5790 2970 5800
rect 3010 5800 3020 5810
rect 3130 5800 3140 5810
rect 3010 5790 3140 5800
rect 3180 5800 3190 5810
rect 3300 5800 3310 5810
rect 3180 5790 3310 5800
rect 3350 5800 3360 5810
rect 3350 5790 3440 5800
rect -60 5770 -50 5790
rect -30 5770 3410 5790
rect 3430 5770 3440 5790
rect -60 5760 30 5770
rect 20 5750 30 5760
rect 70 5760 200 5770
rect 70 5750 80 5760
rect 20 5740 80 5750
rect 190 5750 200 5760
rect 240 5760 370 5770
rect 240 5750 250 5760
rect 190 5740 250 5750
rect 360 5750 370 5760
rect 410 5760 540 5770
rect 410 5750 420 5760
rect 360 5740 420 5750
rect 530 5750 540 5760
rect 580 5760 710 5770
rect 580 5750 590 5760
rect 530 5740 590 5750
rect 700 5750 710 5760
rect 750 5760 880 5770
rect 750 5750 760 5760
rect 700 5740 760 5750
rect 870 5750 880 5760
rect 920 5760 1050 5770
rect 920 5750 930 5760
rect 870 5740 930 5750
rect 1040 5750 1050 5760
rect 1090 5760 1220 5770
rect 1090 5750 1100 5760
rect 1040 5740 1100 5750
rect 1210 5750 1220 5760
rect 1260 5760 1390 5770
rect 1260 5750 1270 5760
rect 1210 5740 1270 5750
rect 1380 5750 1390 5760
rect 1430 5760 1560 5770
rect 1430 5750 1440 5760
rect 1380 5740 1440 5750
rect 1550 5750 1560 5760
rect 1600 5760 1780 5770
rect 1600 5750 1610 5760
rect 1550 5740 1610 5750
rect -310 5690 -270 5700
rect -310 5670 -300 5690
rect -280 5670 -270 5690
rect -310 5640 -270 5670
rect -310 5630 1650 5640
rect -310 5610 -200 5630
rect -160 5610 30 5630
rect 70 5610 200 5630
rect 240 5610 370 5630
rect 410 5610 540 5630
rect 580 5610 710 5630
rect 750 5610 880 5630
rect 920 5610 1050 5630
rect 1090 5610 1220 5630
rect 1260 5610 1390 5630
rect 1430 5610 1560 5630
rect 1600 5610 1650 5630
rect -310 5600 1650 5610
rect -310 1040 -270 5600
rect 1670 5500 1710 5760
rect 1770 5750 1780 5760
rect 1820 5760 1950 5770
rect 1820 5750 1830 5760
rect 1770 5740 1830 5750
rect 1940 5750 1950 5760
rect 1990 5760 2120 5770
rect 1990 5750 2000 5760
rect 1940 5740 2000 5750
rect 2110 5750 2120 5760
rect 2160 5760 2290 5770
rect 2160 5750 2170 5760
rect 2110 5740 2170 5750
rect 2280 5750 2290 5760
rect 2330 5760 2460 5770
rect 2330 5750 2340 5760
rect 2280 5740 2340 5750
rect 2450 5750 2460 5760
rect 2500 5760 2630 5770
rect 2500 5750 2510 5760
rect 2450 5740 2510 5750
rect 2620 5750 2630 5760
rect 2670 5760 2800 5770
rect 2670 5750 2680 5760
rect 2620 5740 2680 5750
rect 2790 5750 2800 5760
rect 2840 5760 2970 5770
rect 2840 5750 2850 5760
rect 2790 5740 2850 5750
rect 2960 5750 2970 5760
rect 3010 5760 3140 5770
rect 3010 5750 3020 5760
rect 2960 5740 3020 5750
rect 3130 5750 3140 5760
rect 3180 5760 3310 5770
rect 3180 5750 3190 5760
rect 3130 5740 3190 5750
rect 3300 5750 3310 5760
rect 3350 5760 3440 5770
rect 3350 5750 3360 5760
rect 3300 5740 3360 5750
rect 3650 5690 3690 5700
rect 3650 5670 3660 5690
rect 3680 5670 3690 5690
rect 3650 5640 3690 5670
rect 1730 5630 3690 5640
rect 1730 5610 1780 5630
rect 1820 5610 1950 5630
rect 1990 5610 2120 5630
rect 2160 5610 2290 5630
rect 2330 5610 2460 5630
rect 2500 5610 2630 5630
rect 2670 5610 2800 5630
rect 2840 5610 2970 5630
rect 3010 5610 3140 5630
rect 3180 5610 3310 5630
rect 3350 5610 3540 5630
rect 3580 5610 3690 5630
rect 1730 5600 3690 5610
rect 20 5490 3360 5500
rect 20 5470 30 5490
rect 70 5470 200 5490
rect 240 5470 370 5490
rect 410 5470 540 5490
rect 580 5470 710 5490
rect 750 5470 880 5490
rect 920 5470 1050 5490
rect 1090 5470 1220 5490
rect 1260 5470 1390 5490
rect 1430 5470 1560 5490
rect 1600 5470 1780 5490
rect 1820 5470 1950 5490
rect 1990 5470 2120 5490
rect 2160 5470 2290 5490
rect 2330 5470 2460 5490
rect 2500 5470 2630 5490
rect 2670 5470 2800 5490
rect 2840 5470 2970 5490
rect 3010 5470 3140 5490
rect 3180 5470 3310 5490
rect 3350 5470 3360 5490
rect 20 5460 3360 5470
rect -210 5090 -110 5100
rect -210 5070 -200 5090
rect -160 5070 -110 5090
rect -210 5060 -110 5070
rect -230 4550 -170 4560
rect -230 4530 -220 4550
rect -180 4530 -170 4550
rect -230 4520 -170 4530
rect -210 4390 -170 4520
rect -210 4370 -200 4390
rect -180 4370 -170 4390
rect -210 4320 -170 4370
rect -150 4400 -110 5060
rect -90 4490 -50 4500
rect -90 4470 -80 4490
rect -60 4470 -50 4490
rect -90 4460 -50 4470
rect -90 4450 1630 4460
rect -90 4430 30 4450
rect 70 4430 200 4450
rect 240 4430 370 4450
rect 410 4430 540 4450
rect 580 4430 710 4450
rect 750 4430 880 4450
rect 920 4430 1050 4450
rect 1090 4430 1220 4450
rect 1260 4430 1390 4450
rect 1430 4430 1560 4450
rect 1600 4430 1630 4450
rect -90 4420 1630 4430
rect 30 4400 70 4420
rect 200 4400 240 4420
rect 370 4400 410 4420
rect 540 4400 580 4420
rect 710 4400 750 4420
rect 880 4400 920 4420
rect 1050 4400 1090 4420
rect 1220 4400 1260 4420
rect 1390 4400 1430 4420
rect 1550 4400 1590 4420
rect -150 4360 -20 4400
rect 30 4390 1590 4400
rect 30 4370 90 4390
rect 110 4370 370 4390
rect 390 4370 650 4390
rect 670 4370 930 4390
rect 950 4370 1210 4390
rect 1230 4370 1590 4390
rect 30 4360 1590 4370
rect -240 4310 -170 4320
rect -240 4270 -230 4310
rect -210 4270 -170 4310
rect -240 4260 -170 4270
rect -210 3870 -170 4260
rect -210 3860 -160 3870
rect -210 3820 -190 3860
rect -170 3820 -160 3860
rect -210 3810 -160 3820
rect -60 3860 -20 4360
rect -60 3820 -50 3860
rect -30 3820 -20 3860
rect -210 3340 -170 3810
rect -60 3790 -20 3820
rect 80 3860 120 4360
rect 80 3820 90 3860
rect 110 3820 120 3860
rect 80 3810 120 3820
rect 220 3860 260 3870
rect 220 3820 230 3860
rect 250 3820 260 3860
rect 220 3790 260 3820
rect 360 3860 400 4360
rect 360 3820 370 3860
rect 390 3820 400 3860
rect 360 3810 400 3820
rect 500 3860 540 3870
rect 500 3820 510 3860
rect 530 3820 540 3860
rect 500 3790 540 3820
rect 640 3860 680 4360
rect 640 3820 650 3860
rect 670 3820 680 3860
rect 640 3810 680 3820
rect 780 3860 820 3870
rect 780 3820 790 3860
rect 810 3820 820 3860
rect 780 3790 820 3820
rect 920 3860 960 4360
rect 920 3820 930 3860
rect 950 3820 960 3860
rect 920 3810 960 3820
rect 1060 3860 1100 3870
rect 1060 3820 1070 3860
rect 1090 3820 1100 3860
rect 1060 3790 1100 3820
rect 1200 3860 1240 4360
rect 1550 4330 1590 4360
rect 1550 4310 1560 4330
rect 1580 4310 1590 4330
rect 1550 4300 1590 4310
rect 1610 4390 1650 4400
rect 1610 4370 1620 4390
rect 1640 4370 1650 4390
rect 1200 3820 1210 3860
rect 1230 3820 1240 3860
rect 1200 3810 1240 3820
rect 1340 3860 1380 3870
rect 1340 3820 1350 3860
rect 1370 3850 1590 3860
rect 1370 3830 1560 3850
rect 1580 3830 1590 3850
rect 1370 3820 1590 3830
rect 1340 3790 1380 3820
rect -60 3750 1380 3790
rect 1610 3485 1650 4370
rect 1610 3415 1620 3485
rect 1640 3415 1650 3485
rect -210 3330 1590 3340
rect -210 3310 1460 3330
rect 1480 3310 1560 3330
rect 1580 3310 1590 3330
rect -210 3300 1590 3310
rect -210 3240 -170 3300
rect -210 3170 -200 3240
rect -180 3170 -170 3240
rect -210 2830 -170 3170
rect -60 2850 1380 2890
rect -210 2820 -160 2830
rect -210 2780 -190 2820
rect -170 2780 -160 2820
rect -210 2770 -160 2780
rect -60 2820 -20 2850
rect -60 2780 -50 2820
rect -30 2780 -20 2820
rect -210 2380 -170 2770
rect -240 2370 -170 2380
rect -240 2330 -230 2370
rect -210 2330 -170 2370
rect -240 2320 -170 2330
rect -210 2270 -170 2320
rect -60 2280 -20 2780
rect 80 2820 120 2830
rect 80 2780 90 2820
rect 110 2780 120 2820
rect 80 2280 120 2780
rect 220 2820 260 2850
rect 220 2780 230 2820
rect 250 2780 260 2820
rect 220 2770 260 2780
rect 360 2820 400 2830
rect 360 2780 370 2820
rect 390 2780 400 2820
rect 360 2280 400 2780
rect 500 2820 540 2850
rect 500 2780 510 2820
rect 530 2780 540 2820
rect 500 2770 540 2780
rect 640 2820 680 2830
rect 640 2780 650 2820
rect 670 2780 680 2820
rect 640 2280 680 2780
rect 780 2820 820 2850
rect 780 2780 790 2820
rect 810 2780 820 2820
rect 780 2770 820 2780
rect 920 2820 960 2830
rect 920 2780 930 2820
rect 950 2780 960 2820
rect 920 2280 960 2780
rect 1060 2820 1100 2850
rect 1060 2780 1070 2820
rect 1090 2780 1100 2820
rect 1060 2770 1100 2780
rect 1200 2820 1240 2830
rect 1200 2780 1210 2820
rect 1230 2780 1240 2820
rect 1200 2280 1240 2780
rect 1340 2820 1380 2850
rect 1340 2780 1350 2820
rect 1370 2810 1590 2820
rect 1370 2790 1560 2810
rect 1580 2790 1590 2810
rect 1370 2780 1590 2790
rect 1340 2770 1380 2780
rect 1550 2330 1590 2340
rect 1550 2310 1560 2330
rect 1580 2310 1590 2330
rect 1550 2280 1590 2310
rect -210 2250 -200 2270
rect -180 2250 -170 2270
rect -210 2120 -170 2250
rect -230 2110 -170 2120
rect -230 2090 -220 2110
rect -180 2090 -170 2110
rect -230 2080 -170 2090
rect -150 2240 -20 2280
rect 30 2270 1590 2280
rect 30 2250 90 2270
rect 110 2250 370 2270
rect 390 2250 650 2270
rect 670 2250 930 2270
rect 950 2250 1210 2270
rect 1230 2250 1590 2270
rect 30 2240 1590 2250
rect 1610 2270 1650 3415
rect 1610 2250 1620 2270
rect 1640 2250 1650 2270
rect 1610 2240 1650 2250
rect -150 1580 -110 2240
rect 30 2220 70 2240
rect 200 2220 240 2240
rect 370 2220 410 2240
rect 540 2220 580 2240
rect 710 2220 750 2240
rect 880 2220 920 2240
rect 1050 2220 1090 2240
rect 1220 2220 1260 2240
rect 1390 2220 1430 2240
rect 1550 2220 1590 2240
rect -90 2210 1630 2220
rect -90 2190 30 2210
rect 70 2190 200 2210
rect 240 2190 370 2210
rect 410 2190 540 2210
rect 580 2190 710 2210
rect 750 2190 880 2210
rect 920 2190 1050 2210
rect 1090 2190 1220 2210
rect 1260 2190 1390 2210
rect 1430 2190 1560 2210
rect 1600 2190 1630 2210
rect -90 2180 1630 2190
rect -90 2170 -50 2180
rect -90 2150 -80 2170
rect -60 2150 -50 2170
rect -90 2140 -50 2150
rect -210 1570 -110 1580
rect -210 1550 -200 1570
rect -160 1550 -110 1570
rect -210 1540 -110 1550
rect 1670 1180 1710 5460
rect 3490 5090 3590 5100
rect 3490 5070 3540 5090
rect 3580 5070 3590 5090
rect 3490 5060 3590 5070
rect 3430 4490 3470 4500
rect 3430 4470 3440 4490
rect 3460 4470 3470 4490
rect 3430 4460 3470 4470
rect 1750 4450 3470 4460
rect 1750 4430 1780 4450
rect 1820 4430 1950 4450
rect 1990 4430 2120 4450
rect 2160 4430 2290 4450
rect 2330 4430 2460 4450
rect 2500 4430 2630 4450
rect 2670 4430 2800 4450
rect 2840 4430 2970 4450
rect 3010 4430 3140 4450
rect 3180 4430 3310 4450
rect 3350 4430 3470 4450
rect 1750 4420 3470 4430
rect 1790 4400 1830 4420
rect 1950 4400 1990 4420
rect 2120 4400 2160 4420
rect 2290 4400 2330 4420
rect 2460 4400 2500 4420
rect 2630 4400 2670 4420
rect 2800 4400 2840 4420
rect 2970 4400 3010 4420
rect 3140 4400 3180 4420
rect 3310 4400 3350 4420
rect 3490 4400 3530 5060
rect 1730 4390 1770 4400
rect 1730 4370 1740 4390
rect 1760 4370 1770 4390
rect 1730 2270 1770 4370
rect 1790 4390 3350 4400
rect 1790 4370 2150 4390
rect 2170 4370 2430 4390
rect 2450 4370 2710 4390
rect 2730 4370 2990 4390
rect 3010 4370 3270 4390
rect 3290 4370 3350 4390
rect 1790 4360 3350 4370
rect 3400 4360 3530 4400
rect 3550 4550 3610 4560
rect 3550 4530 3560 4550
rect 3600 4530 3610 4550
rect 3550 4520 3610 4530
rect 3550 4390 3590 4520
rect 3550 4370 3560 4390
rect 3580 4370 3590 4390
rect 1790 4330 1830 4360
rect 1790 4310 1800 4330
rect 1820 4310 1830 4330
rect 1790 4300 1830 4310
rect 2000 3860 2040 3870
rect 1790 3850 2010 3860
rect 1790 3830 1800 3850
rect 1820 3830 2010 3850
rect 1790 3820 2010 3830
rect 2030 3820 2040 3860
rect 2000 3790 2040 3820
rect 2140 3860 2180 4360
rect 2140 3820 2150 3860
rect 2170 3820 2180 3860
rect 2140 3810 2180 3820
rect 2280 3860 2320 3870
rect 2280 3820 2290 3860
rect 2310 3820 2320 3860
rect 2280 3790 2320 3820
rect 2420 3860 2460 4360
rect 2420 3820 2430 3860
rect 2450 3820 2460 3860
rect 2420 3810 2460 3820
rect 2560 3860 2600 3870
rect 2560 3820 2570 3860
rect 2590 3820 2600 3860
rect 2560 3790 2600 3820
rect 2700 3860 2740 4360
rect 2700 3820 2710 3860
rect 2730 3820 2740 3860
rect 2700 3810 2740 3820
rect 2840 3860 2880 3870
rect 2840 3820 2850 3860
rect 2870 3820 2880 3860
rect 2840 3790 2880 3820
rect 2980 3860 3020 4360
rect 2980 3820 2990 3860
rect 3010 3820 3020 3860
rect 2980 3810 3020 3820
rect 3120 3860 3160 3870
rect 3120 3820 3130 3860
rect 3150 3820 3160 3860
rect 3120 3790 3160 3820
rect 3260 3860 3300 4360
rect 3260 3820 3270 3860
rect 3290 3820 3300 3860
rect 3260 3810 3300 3820
rect 3400 3860 3440 4360
rect 3550 4320 3590 4370
rect 3550 4310 3620 4320
rect 3550 4270 3590 4310
rect 3610 4270 3620 4310
rect 3550 4260 3620 4270
rect 3550 3870 3590 4260
rect 3400 3820 3410 3860
rect 3430 3820 3440 3860
rect 3400 3790 3440 3820
rect 3540 3860 3590 3870
rect 3540 3820 3550 3860
rect 3570 3820 3590 3860
rect 3540 3810 3590 3820
rect 2000 3750 3440 3790
rect 3550 3340 3590 3810
rect 1790 3330 3590 3340
rect 1790 3310 1800 3330
rect 1820 3310 1900 3330
rect 1920 3310 3590 3330
rect 1790 3300 3590 3310
rect 2000 2850 3440 2890
rect 2000 2820 2040 2850
rect 1790 2810 2010 2820
rect 1790 2790 1800 2810
rect 1820 2790 2010 2810
rect 1790 2780 2010 2790
rect 2030 2780 2040 2820
rect 2000 2770 2040 2780
rect 2140 2820 2180 2830
rect 2140 2780 2150 2820
rect 2170 2780 2180 2820
rect 1730 2250 1740 2270
rect 1760 2250 1770 2270
rect 1730 2240 1770 2250
rect 1790 2330 1830 2340
rect 1790 2310 1800 2330
rect 1820 2310 1830 2330
rect 1790 2280 1830 2310
rect 2140 2280 2180 2780
rect 2280 2820 2320 2850
rect 2280 2780 2290 2820
rect 2310 2780 2320 2820
rect 2280 2770 2320 2780
rect 2420 2820 2460 2830
rect 2420 2780 2430 2820
rect 2450 2780 2460 2820
rect 2420 2280 2460 2780
rect 2560 2820 2600 2850
rect 2560 2780 2570 2820
rect 2590 2780 2600 2820
rect 2560 2770 2600 2780
rect 2700 2820 2740 2830
rect 2700 2780 2710 2820
rect 2730 2780 2740 2820
rect 2700 2280 2740 2780
rect 2840 2820 2880 2850
rect 2840 2780 2850 2820
rect 2870 2780 2880 2820
rect 2840 2770 2880 2780
rect 2980 2820 3020 2830
rect 2980 2780 2990 2820
rect 3010 2780 3020 2820
rect 2980 2280 3020 2780
rect 3120 2820 3160 2850
rect 3120 2780 3130 2820
rect 3150 2780 3160 2820
rect 3120 2770 3160 2780
rect 3260 2820 3300 2830
rect 3260 2780 3270 2820
rect 3290 2780 3300 2820
rect 3260 2280 3300 2780
rect 3400 2820 3440 2850
rect 3550 2830 3590 3300
rect 3400 2780 3410 2820
rect 3430 2780 3440 2820
rect 3400 2280 3440 2780
rect 3540 2820 3590 2830
rect 3540 2780 3550 2820
rect 3570 2780 3590 2820
rect 3540 2770 3590 2780
rect 3550 2380 3590 2770
rect 3650 3460 3690 5600
rect 3650 3430 3735 3460
rect 3550 2370 3620 2380
rect 3550 2330 3590 2370
rect 3610 2330 3620 2370
rect 3550 2320 3620 2330
rect 1790 2270 3350 2280
rect 1790 2250 2150 2270
rect 2170 2250 2430 2270
rect 2450 2250 2710 2270
rect 2730 2250 2990 2270
rect 3010 2250 3270 2270
rect 3290 2250 3350 2270
rect 1790 2240 3350 2250
rect 3400 2240 3530 2280
rect 1790 2220 1830 2240
rect 1950 2220 1990 2240
rect 2120 2220 2160 2240
rect 2290 2220 2330 2240
rect 2460 2220 2500 2240
rect 2630 2220 2670 2240
rect 2800 2220 2840 2240
rect 2970 2220 3010 2240
rect 3140 2220 3180 2240
rect 3310 2220 3350 2240
rect 1750 2210 3470 2220
rect 1750 2190 1780 2210
rect 1820 2190 1950 2210
rect 1990 2190 2120 2210
rect 2160 2190 2290 2210
rect 2330 2190 2460 2210
rect 2500 2190 2630 2210
rect 2670 2190 2800 2210
rect 2840 2190 2970 2210
rect 3010 2190 3140 2210
rect 3180 2190 3310 2210
rect 3350 2190 3470 2210
rect 1750 2180 3470 2190
rect 3430 2170 3470 2180
rect 3430 2150 3440 2170
rect 3460 2150 3470 2170
rect 3430 2140 3470 2150
rect 3490 1580 3530 2240
rect 3550 2270 3590 2320
rect 3550 2250 3560 2270
rect 3580 2250 3590 2270
rect 3550 2120 3590 2250
rect 3550 2110 3610 2120
rect 3550 2090 3560 2110
rect 3600 2090 3610 2110
rect 3550 2080 3610 2090
rect 3490 1570 3590 1580
rect 3490 1550 3540 1570
rect 3580 1550 3590 1570
rect 3490 1540 3590 1550
rect 20 1170 3360 1180
rect 20 1150 30 1170
rect 70 1150 200 1170
rect 240 1150 370 1170
rect 410 1150 540 1170
rect 580 1150 710 1170
rect 750 1150 880 1170
rect 920 1150 1050 1170
rect 1090 1150 1220 1170
rect 1260 1150 1390 1170
rect 1430 1150 1560 1170
rect 1600 1150 1780 1170
rect 1820 1150 1950 1170
rect 1990 1150 2120 1170
rect 2160 1150 2290 1170
rect 2330 1150 2460 1170
rect 2500 1150 2630 1170
rect 2670 1150 2800 1170
rect 2840 1150 2970 1170
rect 3010 1150 3140 1170
rect 3180 1150 3310 1170
rect 3350 1150 3360 1170
rect 20 1140 3360 1150
rect -310 1030 1650 1040
rect -310 1010 -200 1030
rect -160 1010 30 1030
rect 70 1010 200 1030
rect 240 1010 370 1030
rect 410 1010 540 1030
rect 580 1010 710 1030
rect 750 1010 880 1030
rect 920 1010 1050 1030
rect 1090 1010 1220 1030
rect 1260 1010 1390 1030
rect 1430 1010 1560 1030
rect 1600 1010 1650 1030
rect -310 1000 1650 1010
rect -310 970 -270 1000
rect -310 950 -300 970
rect -280 950 -270 970
rect -310 940 -270 950
rect 20 890 80 900
rect 20 880 30 890
rect -310 870 30 880
rect 70 880 80 890
rect 190 890 250 900
rect 190 880 200 890
rect 70 870 200 880
rect 240 880 250 890
rect 360 890 420 900
rect 360 880 370 890
rect 240 870 370 880
rect 410 880 420 890
rect 530 890 590 900
rect 530 880 540 890
rect 410 870 540 880
rect 580 880 590 890
rect 700 890 760 900
rect 700 880 710 890
rect 580 870 710 880
rect 750 880 760 890
rect 870 890 930 900
rect 870 880 880 890
rect 750 870 880 880
rect 920 880 930 890
rect 1040 890 1100 900
rect 1040 880 1050 890
rect 920 870 1050 880
rect 1090 880 1100 890
rect 1210 890 1270 900
rect 1210 880 1220 890
rect 1090 870 1220 880
rect 1260 880 1270 890
rect 1380 890 1440 900
rect 1380 880 1390 890
rect 1260 870 1390 880
rect 1430 880 1440 890
rect 1550 890 1610 900
rect 1550 880 1560 890
rect 1430 870 1560 880
rect 1600 880 1610 890
rect 1670 880 1710 1140
rect 3650 1040 3690 3430
rect 1730 1030 3690 1040
rect 1730 1010 1780 1030
rect 1820 1010 1950 1030
rect 1990 1010 2120 1030
rect 2160 1010 2290 1030
rect 2330 1010 2460 1030
rect 2500 1010 2630 1030
rect 2670 1010 2800 1030
rect 2840 1010 2970 1030
rect 3010 1010 3140 1030
rect 3180 1010 3310 1030
rect 3350 1010 3540 1030
rect 3580 1010 3690 1030
rect 1730 1000 3690 1010
rect 3650 970 3690 1000
rect 3650 950 3660 970
rect 3680 950 3690 970
rect 3650 940 3690 950
rect 1770 890 1830 900
rect 1770 880 1780 890
rect 1600 870 1780 880
rect 1820 880 1830 890
rect 1940 890 2000 900
rect 1940 880 1950 890
rect 1820 870 1950 880
rect 1990 880 2000 890
rect 2110 890 2170 900
rect 2110 880 2120 890
rect 1990 870 2120 880
rect 2160 880 2170 890
rect 2280 890 2340 900
rect 2280 880 2290 890
rect 2160 870 2290 880
rect 2330 880 2340 890
rect 2450 890 2510 900
rect 2450 880 2460 890
rect 2330 870 2460 880
rect 2500 880 2510 890
rect 2620 890 2680 900
rect 2620 880 2630 890
rect 2500 870 2630 880
rect 2670 880 2680 890
rect 2790 890 2850 900
rect 2790 880 2800 890
rect 2670 870 2800 880
rect 2840 880 2850 890
rect 2960 890 3020 900
rect 2960 880 2970 890
rect 2840 870 2970 880
rect 3010 880 3020 890
rect 3130 890 3190 900
rect 3130 880 3140 890
rect 3010 870 3140 880
rect 3180 880 3190 890
rect 3300 890 3360 900
rect 3300 880 3310 890
rect 3180 870 3310 880
rect 3350 880 3360 890
rect 3350 870 3690 880
rect -310 850 -50 870
rect -30 850 3410 870
rect 3430 850 3690 870
rect -310 840 30 850
rect 20 830 30 840
rect 70 840 200 850
rect 70 830 80 840
rect 190 830 200 840
rect 240 840 370 850
rect 240 830 250 840
rect 360 830 370 840
rect 410 840 540 850
rect 410 830 420 840
rect 530 830 540 840
rect 580 840 710 850
rect 580 830 590 840
rect 700 830 710 840
rect 750 840 880 850
rect 750 830 760 840
rect 870 830 880 840
rect 920 840 1050 850
rect 920 830 930 840
rect 1040 830 1050 840
rect 1090 840 1220 850
rect 1090 830 1100 840
rect 1210 830 1220 840
rect 1260 840 1390 850
rect 1260 830 1270 840
rect 1380 830 1390 840
rect 1430 840 1560 850
rect 1430 830 1440 840
rect 1550 830 1560 840
rect 1600 840 1780 850
rect 1600 830 1610 840
rect 1770 830 1780 840
rect 1820 840 1950 850
rect 1820 830 1830 840
rect 1940 830 1950 840
rect 1990 840 2120 850
rect 1990 830 2000 840
rect 2110 830 2120 840
rect 2160 840 2290 850
rect 2160 830 2170 840
rect 2280 830 2290 840
rect 2330 840 2460 850
rect 2330 830 2340 840
rect 2450 830 2460 840
rect 2500 840 2630 850
rect 2500 830 2510 840
rect 2620 830 2630 840
rect 2670 840 2800 850
rect 2670 830 2680 840
rect 2790 830 2800 840
rect 2840 840 2970 850
rect 2840 830 2850 840
rect 2960 830 2970 840
rect 3010 840 3140 850
rect 3010 830 3020 840
rect 3130 830 3140 840
rect 3180 840 3310 850
rect 3180 830 3190 840
rect 3300 830 3310 840
rect 3350 840 3690 850
rect 3350 830 3360 840
<< viali >>
rect 1620 3415 1640 3485
rect -200 3170 -180 3240
<< metal1 >>
rect -350 3485 1650 3495
rect -350 3415 1620 3485
rect 1640 3415 1650 3485
rect -350 3405 1650 3415
rect -350 3240 -170 3250
rect -350 3170 -200 3240
rect -180 3170 -170 3240
rect -350 3155 -170 3170
<< labels >>
rlabel locali 3735 3445 3735 3445 3 Vc
port 1 e
rlabel locali 3690 860 3690 860 3 Vp
port 2 e
rlabel metal1 -350 3200 -350 3200 7 Vn
port 4 w
rlabel metal1 -350 3450 -350 3450 7 Vbp
port 3 w
<< end >>
