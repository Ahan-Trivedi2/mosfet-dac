* SPICE3 file created from dac.ext - technology: sky130A


* Top level circuit dac

X0 a_6220_2110# a_6110_n14600# a_6220_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X1 a_2270_n1450# a_n370_n9900# a_2270_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X2 a_3350_n7120# a_n370_n9900# a_3350_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X3 a_1900_3210# a_1790_n14600# a_1900_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X4 a_4060_n7120# a_n370_n9900# a_4060_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X5 a_n370_n5410# a_n370_n5410# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X6 a_110_n350# a_n370_n9900# a_110_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X7 a_n370_n5410# a_n370_n5410# a_3350_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X8 a_3350_n2550# a_n370_n9900# a_2270_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X9 a_n370_n5410# a_n370_n5410# a_4430_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X10 a_4060_n2550# a_n370_n9900# a_3350_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X11 a_4430_n8220# a_n370_n9900# a_4430_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X12 a_5140_n8220# a_n370_n9900# a_5140_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X13 a_5140_4310# a_5030_n14600# a_5140_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X14 a_4060_n10730# a_3950_n14600# a_4060_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X15 a_4430_3210# a_4400_n15030# a_4430_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X16 a_3350_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X17 a_n260_n9320# a_n370_n9900# a_n260_n10730# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X18 a_4430_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X19 a_n370_n5410# a_n370_n5410# a_110_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X20 a_1190_n10420# a_n370_n9900# a_1900_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X21 a_4060_n14030# a_3950_n14600# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X22 a_5140_n11830# a_5030_n14600# a_5140_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X23 a_6220_n10730# a_6560_n15030# a_6590_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X24 a_n370_n5410# a_n370_n5410# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X25 a_n370_n5410# a_n370_n5410# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X26 a_820_n8220# a_n370_n9900# a_820_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X27 a_n260_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X28 a_2270_n9320# a_n370_n9900# a_2270_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X29 a_4430_n350# a_n370_n9900# a_4430_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X30 a_1900_n1450# a_n370_n9900# a_1900_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X31 a_6590_n14030# a_6560_n15030# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X32 a_6220_n12930# a_6110_n14600# a_6220_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X33 a_n370_n5410# a_n370_n5410# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X34 a_5140_n350# a_n370_n9900# a_5140_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X35 a_2270_n10420# a_n370_n9900# a_2980_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X36 a_4430_n10420# a_n370_n9900# a_5510_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X37 a_1900_n12930# a_1790_n14600# a_1900_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X38 a_110_n15130# a_3320_n15030# a_3350_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X39 a_3350_750# a_n370_n9900# a_3350_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X40 a_110_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X41 a_5510_n10420# a_n370_n9900# a_6220_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X42 a_110_3210# a_80_n15030# a_110_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X43 a_820_3210# a_710_n14600# a_820_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X44 a_2980_n1450# a_n370_n9900# a_2980_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X45 a_5510_n1450# a_n370_n9900# a_5510_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X46 a_4060_3210# a_3950_n14600# a_4060_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X47 a_6220_n1450# a_n370_n9900# a_6220_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X48 a_5510_n10420# a_n370_n9900# a_6590_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X49 a_7300_n7120# a_n370_n9900# a_7300_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X50 a_3350_2110# a_3320_n15030# a_2980_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X51 a_820_n350# a_n370_n9900# a_820_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X52 a_n260_n11830# a_n370_n14600# a_n260_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X53 a_110_n15130# a_6560_n15030# a_6590_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X54 a_6590_750# a_n370_n9900# a_6590_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X55 a_820_n10730# a_1160_n15030# a_1190_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X56 a_6590_n1450# a_n370_n9900# a_6590_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X57 a_7300_n2550# a_n370_n9900# a_6590_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X58 a_n260_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X59 a_1190_n14030# a_1160_n15030# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X60 a_2270_n11830# a_2240_n15030# a_2270_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X61 a_6590_2110# a_6560_n15030# a_6220_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X62 a_n370_n5410# a_n370_n5410# a_n260_n6020# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X63 a_5510_n9320# a_n370_n9900# a_5510_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X64 a_2270_4310# a_2240_n15030# a_2270_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X65 a_2980_4310# a_2870_n14600# a_2980_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X66 a_110_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X67 a_3350_n12930# a_3320_n15030# a_3350_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X68 a_n260_n8220# a_n370_n9900# a_n260_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X69 a_110_n12930# a_80_n15030# a_110_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X70 a_n260_n6020# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X71 a_n370_n5410# a_n370_n5410# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X72 a_4060_n10730# a_4400_n15030# a_4430_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X73 a_820_n9320# a_n370_n9900# a_820_n10730# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X74 a_110_n15130# a_n370_n9900# a_7300_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X75 a_n370_n5410# a_n370_n5410# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X76 a_n260_n350# a_n370_n9900# a_n260_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X77 a_4430_n14030# a_4400_n15030# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X78 a_5510_n11830# a_5480_n15030# a_5510_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X79 a_1190_3210# a_1160_n15030# a_1190_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X80 a_1190_n7120# a_n370_n9900# a_1190_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X81 a_2980_n10730# a_2870_n14600# a_2980_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X82 a_n370_n5410# a_n370_n5410# a_1190_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X83 a_110_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X84 a_n260_3210# a_n370_n14600# a_n260_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X85 a_2980_n14030# a_2870_n14600# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X86 a_n370_n5410# a_n370_n5410# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X87 a_1190_n2550# a_n370_n9900# a_110_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X88 a_2270_n8220# a_n370_n9900# a_2270_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X89 a_110_n7120# a_n370_n9900# a_110_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X90 a_820_n11830# a_710_n14600# a_820_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X91 a_6220_4310# a_6110_n14600# a_6220_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X92 a_5510_3210# a_5480_n15030# a_5510_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X93 a_1190_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X94 a_n260_n15130# a_1790_n14600# a_1900_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X95 a_1900_750# a_n370_n9900# a_1900_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X96 a_110_n2550# a_n370_n9900# a_n260_n6020# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X97 a_n260_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X98 a_2270_n350# a_n370_n9900# a_2270_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X99 a_2270_n10420# a_n370_n9900# a_3350_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X100 a_1900_2110# a_1790_n14600# a_1900_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X101 a_3350_n10420# a_n370_n9900# a_4060_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X102 a_6220_n9320# a_n370_n9900# a_6220_n10730# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X103 a_n370_n5410# a_n370_n5410# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X104 a_110_n15130# a_4400_n15030# a_4430_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X105 a_n370_n5410# a_n370_n5410# a_1190_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X106 a_4060_n12930# a_3950_n14600# a_4060_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X107 a_1900_n9320# a_n370_n9900# a_1900_n10730# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X108 a_4430_750# a_n370_n9900# a_4430_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X109 a_3350_n1450# a_n370_n9900# a_3350_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X110 a_4060_n1450# a_n370_n9900# a_4060_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X111 a_4430_n7120# a_n370_n9900# a_4430_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X112 a_1900_n8220# a_n370_n9900# a_1900_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X113 a_5140_n7120# a_n370_n9900# a_5140_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X114 a_6590_n12930# a_6560_n15030# a_6590_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X115 a_5140_3210# a_5030_n14600# a_5140_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X116 a_n370_n5410# a_n370_n5410# a_2270_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X117 a_n370_n5410# a_n370_n5410# a_4430_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X118 a_n370_n5410# a_n370_n5410# a_5510_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X119 a_4430_2110# a_4400_n15030# a_4060_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X120 a_4430_n2550# a_n370_n9900# a_3350_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X121 a_1190_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X122 a_5140_n2550# a_n370_n9900# a_4430_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X123 a_5140_n10730# a_5030_n14600# a_5140_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X124 a_5510_n8220# a_n370_n9900# a_5510_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X125 a_2980_n8220# a_n370_n9900# a_2980_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X126 a_6220_n8220# a_n370_n9900# a_6220_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X127 a_110_n15130# a_80_n15030# a_110_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X128 a_n260_n15130# a_710_n14600# a_820_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X129 a_110_750# a_n370_n9900# a_110_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X130 a_820_750# a_n370_n9900# a_820_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X131 a_n370_n5410# a_n370_n5410# a_5510_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X132 a_820_n7120# a_n370_n9900# a_820_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X133 a_1900_n350# a_n370_n9900# a_1900_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X134 a_2270_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X135 a_4430_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X136 a_5140_n14030# a_5030_n14600# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X137 a_6220_n11830# a_6110_n14600# a_6220_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X138 a_n260_n15130# a_3950_n14600# a_4060_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X139 a_4060_750# a_n370_n9900# a_4060_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X140 a_5510_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X141 a_1900_n11830# a_1790_n14600# a_1900_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X142 a_6590_n8220# a_n370_n9900# a_6590_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X143 a_3350_4310# a_3320_n15030# a_3350_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X144 a_820_n2550# a_n370_n9900# a_110_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X145 a_n260_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X146 a_3350_n9320# a_n370_n9900# a_3350_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X147 a_110_2110# a_80_n15030# a_n260_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X148 a_820_2110# a_710_n14600# a_820_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X149 a_n260_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X150 a_1190_n12930# a_1160_n15030# a_1190_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X151 a_2980_n350# a_n370_n9900# a_2980_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X152 a_5510_n350# a_n370_n9900# a_5510_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X153 a_5510_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X154 a_4060_2110# a_3950_n14600# a_4060_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X155 a_6220_n350# a_n370_n9900# a_6220_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X156 a_110_n9320# a_n370_n9900# a_110_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X157 a_6590_n10420# a_n370_n9900# a_7300_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X158 a_n260_n10730# a_n370_n14600# a_n260_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X159 a_6590_4310# a_6560_n15030# a_6590_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X160 a_n370_n5410# a_n370_n5410# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X161 a_n370_n5410# a_n370_n5410# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X162 a_6590_n350# a_n370_n9900# a_6590_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X163 a_7300_n1450# a_n370_n9900# a_7300_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X164 a_n260_n14030# a_n370_n14600# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X165 a_1900_n10730# a_2240_n15030# a_2270_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X166 a_2270_3210# a_2240_n15030# a_2270_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X167 a_2980_3210# a_2870_n14600# a_2980_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X168 a_2270_n14030# a_2240_n15030# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X169 a_3350_n11830# a_3320_n15030# a_3350_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X170 a_n260_n7120# a_n370_n9900# a_n260_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X171 a_110_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X172 a_4430_n12930# a_4400_n15030# a_4430_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X173 a_110_n11830# a_80_n15030# a_110_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X174 a_n260_n2550# a_n370_n9900# a_n260_n6020# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X175 a_110_n15130# a_1160_n15030# a_1190_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X176 a_1190_750# a_n370_n9900# a_1190_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X177 a_110_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X178 a_2980_n12930# a_2870_n14600# a_2980_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X179 a_n260_n15130# a_n370_n14600# a_n260_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X180 a_n260_750# a_n370_n9900# a_n260_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X181 a_5140_n10730# a_5480_n15030# a_5510_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X182 a_1190_2110# a_1160_n15030# a_820_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X183 a_110_n10420# a_n370_n9900# a_1190_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X184 a_5510_n14030# a_5480_n15030# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X185 a_n260_2110# a_n370_n14600# a_n260_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X186 a_n370_n5410# a_n370_n5410# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X187 a_110_n15130# a_5480_n15030# a_5510_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X188 a_1190_n1450# a_n370_n9900# a_1190_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X189 a_4060_n9320# a_n370_n9900# a_4060_n10730# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X190 a_5510_750# a_n370_n9900# a_5510_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X191 a_2270_n7120# a_n370_n9900# a_2270_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X192 a_n370_n5410# a_n370_n5410# a_2270_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X193 a_6590_n9320# a_n370_n9900# a_6590_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X194 a_n370_n5410# a_n370_n5410# a_3350_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X195 a_n260_n6020# a_n370_n9900# a_110_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X196 a_820_n10730# a_710_n14600# a_820_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X197 a_6220_3210# a_6110_n14600# a_6220_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X198 a_5510_2110# a_5480_n15030# a_5140_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X199 a_2270_n2550# a_n370_n9900# a_1190_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X200 a_3350_n8220# a_n370_n9900# a_3350_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X201 a_1900_4310# a_1790_n14600# a_1900_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X202 a_820_n14030# a_710_n14600# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X203 a_4060_n8220# a_n370_n9900# a_4060_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X204 a_110_n1450# a_n370_n9900# a_110_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X205 a_2270_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X206 a_3350_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X207 a_n260_n15130# a_5030_n14600# a_5140_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X208 a_5140_750# a_n370_n9900# a_5140_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X209 a_4060_n11830# a_3950_n14600# a_4060_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X210 a_4430_4310# a_4400_n15030# a_4430_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X211 a_7300_n9320# a_n370_n9900# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X212 a_3350_n350# a_n370_n9900# a_3350_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X213 a_4060_n350# a_n370_n9900# a_4060_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X214 a_3350_n10420# a_n370_n9900# a_4430_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X215 a_1900_n7120# a_n370_n9900# a_1900_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X216 a_n260_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X217 a_5140_n12930# a_5030_n14600# a_5140_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X218 a_1190_n9320# a_n370_n9900# a_1190_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X219 a_4430_n10420# a_n370_n9900# a_5140_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X220 a_6590_n11830# a_6560_n15030# a_6590_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X221 a_5140_2110# a_5030_n14600# a_5140_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X222 a_4430_n1450# a_n370_n9900# a_4430_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X223 a_1900_n2550# a_n370_n9900# a_1190_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X224 a_110_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X225 a_5140_n1450# a_n370_n9900# a_5140_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X226 a_2980_n7120# a_n370_n9900# a_2980_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X227 a_5510_n7120# a_n370_n9900# a_5510_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X228 a_n370_n5410# a_n370_n5410# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X229 a_6220_n7120# a_n370_n9900# a_6220_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X230 a_110_4310# a_80_n15030# a_110_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X231 a_820_4310# a_710_n14600# a_820_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X232 a_n370_n5410# a_n370_n5410# a_6590_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X233 a_110_n10420# a_n370_n9900# a_820_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X234 a_2980_n2550# a_n370_n9900# a_2270_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X235 a_5510_n2550# a_n370_n9900# a_4430_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X236 a_6220_n10730# a_6110_n14600# a_6220_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X237 a_4060_4310# a_3950_n14600# a_4060_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X238 a_6220_n2550# a_n370_n9900# a_5510_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X239 a_6590_n7120# a_n370_n9900# a_6590_n8220# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X240 a_1900_n10730# a_1790_n14600# a_1900_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X241 a_7300_n8220# a_n370_n9900# a_7300_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X242 a_3350_3210# a_3320_n15030# a_3350_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X243 a_820_n1450# a_n370_n9900# a_820_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X244 a_6220_n14030# a_6110_n14600# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X245 a_n260_n12930# a_n370_n14600# a_n260_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X246 a_n370_n5410# a_n370_n5410# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X247 a_1900_n14030# a_1790_n14600# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X248 a_1190_n11830# a_1160_n15030# a_1190_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X249 a_6590_n2550# a_n370_n9900# a_5510_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X250 a_6590_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X251 a_4430_n9320# a_n370_n9900# a_4430_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X252 a_110_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X253 a_2270_n12930# a_2240_n15030# a_2270_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X254 a_6590_3210# a_6560_n15030# a_6590_2110# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X255 a_2980_n9320# a_n370_n9900# a_2980_n10730# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X256 a_110_n15130# a_2240_n15030# a_2270_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X257 a_n260_n15130# a_2870_n14600# a_2980_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X258 a_2270_750# a_n370_n9900# a_2270_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X259 a_2980_750# a_n370_n9900# a_2980_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X260 a_7300_n350# a_n370_n9900# a_7300_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X261 a_2270_2110# a_2240_n15030# a_1900_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X262 a_2980_2110# a_2870_n14600# a_2980_750# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X263 a_2980_n10730# a_3320_n15030# a_3350_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X264 a_n260_n6020# a_n370_n9900# a_n260_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X265 a_3350_n14030# a_3320_n15030# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X266 a_4430_n11830# a_4400_n15030# a_4430_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X267 a_n370_n5410# a_n370_n5410# a_110_n10420# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X268 a_110_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X269 a_n260_n10730# a_80_n15030# a_110_n11830# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X270 a_n260_n1450# a_n370_n9900# a_n260_n2550# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X271 a_5510_n12930# a_5480_n15030# a_5510_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X272 a_1190_4310# a_1160_n15030# a_1190_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X273 a_1190_n8220# a_n370_n9900# a_1190_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X274 a_110_n14030# a_80_n15030# a_110_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X275 a_2980_n11830# a_2870_n14600# a_2980_n12930# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X276 a_n260_4310# a_n370_n14600# a_n260_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X277 a_n260_n15130# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X278 a_110_750# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X279 a_n370_n5410# a_n370_n5410# a_n260_n6020# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X280 a_110_n8220# a_n370_n9900# a_110_n9320# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X281 a_820_n12930# a_710_n14600# a_820_n14030# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X282 a_n260_n15130# a_6110_n14600# a_6220_4310# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X283 a_5510_4310# a_5480_n15030# a_5510_3210# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X284 a_6220_750# a_n370_n9900# a_6220_n350# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X285 a_1190_n350# a_n370_n9900# a_1190_n1450# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X286 a_n370_n5410# a_n370_n5410# a_n260_n15130# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X287 a_n260_n6020# a_n370_n5410# a_n370_n5410# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X288 a_1190_n10420# a_n370_n9900# a_2270_n7120# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X289 a_5140_n9320# a_n370_n9900# a_5140_n10730# a_n370_n5410# sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
.end

