magic
tech sky130A
timestamp 1762139857
<< locali >>
rect 6865 7905 6945 7910
rect 6865 7885 6870 7905
rect 6940 7885 6945 7905
rect 6865 7875 6945 7885
rect 6800 5315 6915 5325
rect 6800 5295 6810 5315
rect 6880 5295 6915 5315
rect 6800 5285 6915 5295
rect 2040 830 2080 840
rect 2040 760 2050 830
rect 2070 760 2080 830
rect 2040 750 2080 760
rect 2195 830 2235 840
rect 2195 760 2205 830
rect 2225 760 2235 830
rect 2195 40 2235 760
rect 2040 20 2235 40
<< viali >>
rect 6870 7885 6940 7905
rect 2870 5295 2940 5315
rect 6810 5295 6880 5315
rect 2050 760 2070 830
rect 2205 760 2225 830
rect 2840 25 2910 45
<< metal1 >>
rect 2040 7850 4380 7940
rect 4760 7850 6745 7940
rect 6855 7905 6965 7910
rect 6855 7885 6870 7905
rect 6940 7885 6965 7905
rect 6855 7875 6965 7885
rect 2040 830 2080 7850
rect 2770 5520 2805 7695
rect 2970 7595 6395 7695
rect 6300 6680 6395 7595
rect 6705 7275 6745 7850
rect 6705 6950 6750 7275
rect 6710 6865 6750 6950
rect 6930 6910 6965 7875
rect 6930 6885 7465 6910
rect 6705 6855 7400 6865
rect 6705 6815 7200 6855
rect 6710 6810 6750 6815
rect 7185 6785 7200 6815
rect 7230 6815 7400 6855
rect 7230 6785 7245 6815
rect 7510 6800 7540 6875
rect 7185 6780 7245 6785
rect 7500 6785 7540 6800
rect 7500 6715 7505 6785
rect 7535 6715 7540 6785
rect 7500 6705 7540 6715
rect 6300 6590 7890 6680
rect 7555 5925 7635 6590
rect 7555 5825 7575 5925
rect 7615 5825 7635 5925
rect 7555 5810 7635 5825
rect 6980 5675 7745 5715
rect 8390 5675 8415 5680
rect 2765 5510 2815 5520
rect 2765 5440 2775 5510
rect 2805 5440 2815 5510
rect 2765 5430 2815 5440
rect 2410 5325 2735 5330
rect 6980 5325 7035 5675
rect 2410 5315 2950 5325
rect 2410 5295 2870 5315
rect 2940 5295 2950 5315
rect 2410 5285 2950 5295
rect 6800 5315 7035 5325
rect 6800 5295 6810 5315
rect 6880 5295 7035 5315
rect 6800 5285 7035 5295
rect 2410 2785 2485 5285
rect 8390 4955 8420 5675
rect 7365 3620 7525 3645
rect 7365 3550 7480 3620
rect 7510 3550 7525 3620
rect 7365 3530 7525 3550
rect 7365 3350 7410 3530
rect 7185 3340 7245 3350
rect 7185 3270 7200 3340
rect 7230 3300 7245 3340
rect 7365 3325 7455 3350
rect 7230 3270 7455 3300
rect 7185 3255 7455 3270
rect 2410 2715 2430 2785
rect 2460 2715 2485 2785
rect 2410 2705 2485 2715
rect 2040 760 2050 830
rect 2070 760 2080 830
rect 2040 750 2080 760
rect 2190 2185 2875 2285
rect 2190 830 2255 2185
rect 2190 760 2205 830
rect 2225 760 2255 830
rect 2190 745 2255 760
rect 2415 2125 2800 2150
rect 2415 2055 2430 2125
rect 2460 2055 2800 2125
rect 2415 2050 2800 2055
rect 2415 655 2480 2050
rect 2040 560 2480 655
rect 2755 80 2820 90
rect 2755 20 2775 80
rect 2040 10 2775 20
rect 2805 60 2820 80
rect 2805 45 2920 60
rect 2805 25 2840 45
rect 2910 25 2920 45
rect 2805 10 2920 25
rect 2040 0 2920 10
<< via1 >>
rect 7200 6785 7230 6855
rect 7505 6715 7535 6785
rect 7575 5825 7615 5925
rect 2775 5440 2805 5510
rect 7480 3550 7510 3620
rect 7200 3270 7230 3340
rect 7945 3040 7975 3110
rect 2430 2715 2460 2785
rect 2430 2055 2460 2125
rect 2775 10 2805 80
<< metal2 >>
rect 7185 6855 7245 6865
rect 7185 6785 7200 6855
rect 7230 6785 7245 6855
rect 2765 5510 2815 5520
rect 2765 5440 2775 5510
rect 2805 5440 2815 5510
rect 2420 2785 2470 2805
rect 2420 2715 2430 2785
rect 2460 2715 2470 2785
rect 2420 2125 2470 2715
rect 2420 2055 2430 2125
rect 2460 2055 2470 2125
rect 2420 2045 2470 2055
rect 2765 80 2815 5440
rect 7185 3340 7245 6785
rect 7500 6785 7540 6800
rect 7500 6715 7505 6785
rect 7535 6715 7540 6785
rect 7500 3640 7540 6715
rect 7555 5925 7635 5970
rect 7555 5825 7575 5925
rect 7615 5825 7635 5925
rect 7555 5810 7635 5825
rect 7560 4460 7635 5810
rect 7560 4390 7645 4460
rect 7560 4385 7940 4390
rect 7560 4280 7995 4385
rect 7465 3620 7540 3640
rect 7465 3550 7480 3620
rect 7510 3550 7540 3620
rect 7465 3535 7540 3550
rect 7185 3270 7200 3340
rect 7230 3270 7245 3340
rect 7185 3260 7245 3270
rect 7920 3110 7995 4280
rect 7920 3040 7945 3110
rect 7975 3040 7995 3110
rect 7920 3010 7995 3040
rect 2765 10 2775 80
rect 2805 10 2815 80
rect 2765 0 2815 10
use bbg  bbg_0
timestamp 1762117721
transform 1 0 220 0 1 560
box -220 -560 1820 210
use ccm  ccm_0
timestamp 1762061669
transform 1 0 9265 0 1 25
box -1810 -10 2910 1120
use fvf  fvf_0
timestamp 1762117721
transform 0 1 7910 -1 0 8390
box -150 -510 3125 510
use fvf  fvf_1
timestamp 1762117721
transform 0 1 7960 -1 0 4830
box -150 -510 3125 510
use ncbc  ncbc_0
timestamp 1762137910
transform 1 0 3155 0 1 4445
box -350 810 3735 5830
use pcbc  pcbc_0
timestamp 1762135317
transform 1 0 -1317 0 1 -2702
box 4115 2710 8150 7690
<< end >>
