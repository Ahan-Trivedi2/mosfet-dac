magic
tech sky130A
timestamp 1762032340
<< nwell >>
rect -310 2710 3690 5110
rect -310 -90 3690 2310
<< nmos >>
rect -160 2560 -60 2660
rect -20 2560 80 2660
rect 120 2560 220 2660
rect 260 2560 360 2660
rect 400 2560 500 2660
rect 540 2560 640 2660
rect 680 2560 780 2660
rect 820 2560 920 2660
rect 960 2560 1060 2660
rect 1100 2560 1200 2660
rect 1240 2560 1340 2660
rect 2040 2560 2140 2660
rect 2180 2560 2280 2660
rect 2320 2560 2420 2660
rect 2460 2560 2560 2660
rect 2600 2560 2700 2660
rect 2740 2560 2840 2660
rect 2880 2560 2980 2660
rect 3020 2560 3120 2660
rect 3160 2560 3260 2660
rect 3300 2560 3400 2660
rect 3440 2560 3540 2660
rect -160 2360 -60 2460
rect -20 2360 80 2460
rect 120 2360 220 2460
rect 260 2360 360 2460
rect 400 2360 500 2460
rect 540 2360 640 2460
rect 680 2360 780 2460
rect 820 2360 920 2460
rect 960 2360 1060 2460
rect 1100 2360 1200 2460
rect 1240 2360 1340 2460
rect 2040 2360 2140 2460
rect 2180 2360 2280 2460
rect 2320 2360 2420 2460
rect 2460 2360 2560 2460
rect 2600 2360 2700 2460
rect 2740 2360 2840 2460
rect 2880 2360 2980 2460
rect 3020 2360 3120 2460
rect 3160 2360 3260 2460
rect 3300 2360 3400 2460
rect 3440 2360 3540 2460
<< pmos >>
rect 0 4020 100 5020
rect 170 4020 270 5020
rect 340 4020 440 5020
rect 510 4020 610 5020
rect 680 4020 780 5020
rect 850 4020 950 5020
rect 1020 4020 1120 5020
rect 1190 4020 1290 5020
rect 1360 4020 1460 5020
rect 1530 4020 1630 5020
rect 1750 4020 1850 5020
rect 1920 4020 2020 5020
rect 2090 4020 2190 5020
rect 2260 4020 2360 5020
rect 2430 4020 2530 5020
rect 2600 4020 2700 5020
rect 2770 4020 2870 5020
rect 2940 4020 3040 5020
rect 3110 4020 3210 5020
rect 3280 4020 3380 5020
rect -280 3480 -80 3980
rect -280 2940 -80 3440
rect 0 2980 100 3980
rect 170 2980 270 3980
rect 340 2980 440 3980
rect 510 2980 610 3980
rect 680 2980 780 3980
rect 850 2980 950 3980
rect 1020 2980 1120 3980
rect 1190 2980 1290 3980
rect 1360 2980 1460 3980
rect 1530 2980 1630 3980
rect 0 2770 100 2870
rect 170 2770 270 2870
rect 340 2770 440 2870
rect 510 2770 610 2870
rect 680 2770 780 2870
rect 850 2770 950 2870
rect 1020 2770 1120 2870
rect 1190 2770 1290 2870
rect 1360 2770 1460 2870
rect 1530 2770 1630 2870
rect 1750 2980 1850 3980
rect 1920 2980 2020 3980
rect 2090 2980 2190 3980
rect 2260 2980 2360 3980
rect 2430 2980 2530 3980
rect 2600 2980 2700 3980
rect 2770 2980 2870 3980
rect 2940 2980 3040 3980
rect 3110 2980 3210 3980
rect 3280 2980 3380 3980
rect 3460 3480 3660 3980
rect 3460 2940 3660 3440
rect 1750 2770 1850 2870
rect 1920 2770 2020 2870
rect 2090 2770 2190 2870
rect 2260 2770 2360 2870
rect 2430 2770 2530 2870
rect 2600 2770 2700 2870
rect 2770 2770 2870 2870
rect 2940 2770 3040 2870
rect 3110 2770 3210 2870
rect 3280 2770 3380 2870
rect 0 2150 100 2250
rect 170 2150 270 2250
rect 340 2150 440 2250
rect 510 2150 610 2250
rect 680 2150 780 2250
rect 850 2150 950 2250
rect 1020 2150 1120 2250
rect 1190 2150 1290 2250
rect 1360 2150 1460 2250
rect 1530 2150 1630 2250
rect -280 1580 -80 2080
rect -280 1040 -80 1540
rect 0 1040 100 2040
rect 170 1040 270 2040
rect 340 1040 440 2040
rect 510 1040 610 2040
rect 680 1040 780 2040
rect 850 1040 950 2040
rect 1020 1040 1120 2040
rect 1190 1040 1290 2040
rect 1360 1040 1460 2040
rect 1530 1040 1630 2040
rect 1750 2150 1850 2250
rect 1920 2150 2020 2250
rect 2090 2150 2190 2250
rect 2260 2150 2360 2250
rect 2430 2150 2530 2250
rect 2600 2150 2700 2250
rect 2770 2150 2870 2250
rect 2940 2150 3040 2250
rect 3110 2150 3210 2250
rect 3280 2150 3380 2250
rect 1750 1040 1850 2040
rect 1920 1040 2020 2040
rect 2090 1040 2190 2040
rect 2260 1040 2360 2040
rect 2430 1040 2530 2040
rect 2600 1040 2700 2040
rect 2770 1040 2870 2040
rect 2940 1040 3040 2040
rect 3110 1040 3210 2040
rect 3280 1040 3380 2040
rect 3460 1580 3660 2080
rect 3460 1040 3660 1540
rect 0 0 100 1000
rect 170 0 270 1000
rect 340 0 440 1000
rect 510 0 610 1000
rect 680 0 780 1000
rect 850 0 950 1000
rect 1020 0 1120 1000
rect 1190 0 1290 1000
rect 1360 0 1460 1000
rect 1530 0 1630 1000
rect 1750 0 1850 1000
rect 1920 0 2020 1000
rect 2090 0 2190 1000
rect 2260 0 2360 1000
rect 2430 0 2530 1000
rect 2600 0 2700 1000
rect 2770 0 2870 1000
rect 2940 0 3040 1000
rect 3110 0 3210 1000
rect 3280 0 3380 1000
<< ndiff >>
rect 1550 2660 1590 2670
rect 1790 2660 1830 2670
rect -240 2650 -160 2660
rect -200 2630 -160 2650
rect -200 2590 -190 2630
rect -170 2590 -160 2630
rect -200 2560 -160 2590
rect -60 2630 -20 2660
rect -60 2590 -50 2630
rect -30 2590 -20 2630
rect -60 2560 -20 2590
rect 80 2630 120 2660
rect 80 2590 90 2630
rect 110 2590 120 2630
rect 80 2560 120 2590
rect 220 2630 260 2660
rect 220 2590 230 2630
rect 250 2590 260 2630
rect 220 2560 260 2590
rect 360 2630 400 2660
rect 360 2590 370 2630
rect 390 2590 400 2630
rect 360 2560 400 2590
rect 500 2630 540 2660
rect 500 2590 510 2630
rect 530 2590 540 2630
rect 500 2560 540 2590
rect 640 2630 680 2660
rect 640 2590 650 2630
rect 670 2590 680 2630
rect 640 2560 680 2590
rect 780 2630 820 2660
rect 780 2590 790 2630
rect 810 2590 820 2630
rect 780 2560 820 2590
rect 920 2630 960 2660
rect 920 2590 930 2630
rect 950 2590 960 2630
rect 920 2560 960 2590
rect 1060 2630 1100 2660
rect 1060 2590 1070 2630
rect 1090 2590 1100 2630
rect 1060 2560 1100 2590
rect 1200 2630 1240 2660
rect 1200 2590 1210 2630
rect 1230 2590 1240 2630
rect 1200 2560 1240 2590
rect 1340 2630 1380 2660
rect 1550 2640 1560 2660
rect 1580 2640 1800 2660
rect 1820 2640 1830 2660
rect 1550 2630 1830 2640
rect 2000 2630 2040 2660
rect 1340 2590 1350 2630
rect 1370 2590 1380 2630
rect 1340 2560 1380 2590
rect 1550 2590 1830 2600
rect 1550 2570 1560 2590
rect 1580 2570 1800 2590
rect 1820 2570 1830 2590
rect 1550 2560 1830 2570
rect 2000 2590 2010 2630
rect 2030 2590 2040 2630
rect 2000 2560 2040 2590
rect 2140 2630 2180 2660
rect 2140 2590 2150 2630
rect 2170 2590 2180 2630
rect 2140 2560 2180 2590
rect 2280 2630 2320 2660
rect 2280 2590 2290 2630
rect 2310 2590 2320 2630
rect 2280 2560 2320 2590
rect 2420 2630 2460 2660
rect 2420 2590 2430 2630
rect 2450 2590 2460 2630
rect 2420 2560 2460 2590
rect 2560 2630 2600 2660
rect 2560 2590 2570 2630
rect 2590 2590 2600 2630
rect 2560 2560 2600 2590
rect 2700 2630 2740 2660
rect 2700 2590 2710 2630
rect 2730 2590 2740 2630
rect 2700 2560 2740 2590
rect 2840 2630 2880 2660
rect 2840 2590 2850 2630
rect 2870 2590 2880 2630
rect 2840 2560 2880 2590
rect 2980 2630 3020 2660
rect 2980 2590 2990 2630
rect 3010 2590 3020 2630
rect 2980 2560 3020 2590
rect 3120 2630 3160 2660
rect 3120 2590 3130 2630
rect 3150 2590 3160 2630
rect 3120 2560 3160 2590
rect 3260 2630 3300 2660
rect 3260 2590 3270 2630
rect 3290 2590 3300 2630
rect 3260 2560 3300 2590
rect 3400 2630 3440 2660
rect 3400 2590 3410 2630
rect 3430 2590 3440 2630
rect 3400 2560 3440 2590
rect 3540 2650 3620 2660
rect 3540 2630 3580 2650
rect 3540 2590 3550 2630
rect 3570 2590 3580 2630
rect 3540 2560 3580 2590
rect 1210 2460 1230 2560
rect 1350 2460 1370 2560
rect 1550 2520 1830 2530
rect 1550 2500 1560 2520
rect 1580 2500 1800 2520
rect 1820 2500 1830 2520
rect 1550 2490 1830 2500
rect 2010 2460 2030 2560
rect 2150 2460 2170 2560
rect -200 2430 -160 2460
rect -200 2390 -190 2430
rect -170 2390 -160 2430
rect -200 2370 -160 2390
rect -240 2360 -160 2370
rect -60 2430 -20 2460
rect -60 2390 -50 2430
rect -30 2390 -20 2430
rect -60 2360 -20 2390
rect 80 2430 120 2460
rect 80 2390 90 2430
rect 110 2390 120 2430
rect 80 2360 120 2390
rect 220 2430 260 2460
rect 220 2390 230 2430
rect 250 2390 260 2430
rect 220 2360 260 2390
rect 360 2430 400 2460
rect 360 2390 370 2430
rect 390 2390 400 2430
rect 360 2360 400 2390
rect 500 2430 540 2460
rect 500 2390 510 2430
rect 530 2390 540 2430
rect 500 2360 540 2390
rect 640 2430 680 2460
rect 640 2390 650 2430
rect 670 2390 680 2430
rect 640 2360 680 2390
rect 780 2430 820 2460
rect 780 2390 790 2430
rect 810 2390 820 2430
rect 780 2360 820 2390
rect 920 2430 960 2460
rect 920 2390 930 2430
rect 950 2390 960 2430
rect 920 2360 960 2390
rect 1060 2430 1100 2460
rect 1060 2390 1070 2430
rect 1090 2390 1100 2430
rect 1060 2360 1100 2390
rect 1200 2430 1240 2460
rect 1200 2390 1210 2430
rect 1230 2390 1240 2430
rect 1200 2360 1240 2390
rect 1340 2430 1380 2460
rect 1340 2390 1350 2430
rect 1370 2390 1380 2430
rect 1550 2450 1830 2460
rect 1550 2430 1560 2450
rect 1580 2430 1800 2450
rect 1820 2430 1830 2450
rect 1550 2420 1830 2430
rect 2000 2430 2040 2460
rect 2000 2390 2010 2430
rect 2030 2390 2040 2430
rect 1340 2360 1380 2390
rect 1550 2380 1830 2390
rect 1550 2360 1560 2380
rect 1580 2360 1800 2380
rect 1820 2360 1830 2380
rect 2000 2360 2040 2390
rect 2140 2430 2180 2460
rect 2140 2390 2150 2430
rect 2170 2390 2180 2430
rect 2140 2360 2180 2390
rect 2280 2430 2320 2460
rect 2280 2390 2290 2430
rect 2310 2390 2320 2430
rect 2280 2360 2320 2390
rect 2420 2430 2460 2460
rect 2420 2390 2430 2430
rect 2450 2390 2460 2430
rect 2420 2360 2460 2390
rect 2560 2430 2600 2460
rect 2560 2390 2570 2430
rect 2590 2390 2600 2430
rect 2560 2360 2600 2390
rect 2700 2430 2740 2460
rect 2700 2390 2710 2430
rect 2730 2390 2740 2430
rect 2700 2360 2740 2390
rect 2840 2430 2880 2460
rect 2840 2390 2850 2430
rect 2870 2390 2880 2430
rect 2840 2360 2880 2390
rect 2980 2430 3020 2460
rect 2980 2390 2990 2430
rect 3010 2390 3020 2430
rect 2980 2360 3020 2390
rect 3120 2430 3160 2460
rect 3120 2390 3130 2430
rect 3150 2390 3160 2430
rect 3120 2360 3160 2390
rect 3260 2430 3300 2460
rect 3260 2390 3270 2430
rect 3290 2390 3300 2430
rect 3260 2360 3300 2390
rect 3400 2430 3440 2460
rect 3400 2390 3410 2430
rect 3430 2390 3440 2430
rect 3400 2360 3440 2390
rect 3540 2430 3580 2460
rect 3540 2390 3550 2430
rect 3570 2390 3580 2430
rect 3540 2370 3580 2390
rect 3540 2360 3620 2370
rect 1550 2350 1590 2360
rect 1790 2350 1830 2360
<< pdiff >>
rect 0 5050 100 5060
rect 0 5030 30 5050
rect 70 5030 100 5050
rect 0 5020 100 5030
rect 170 5050 270 5060
rect 170 5030 200 5050
rect 240 5030 270 5050
rect 170 5020 270 5030
rect 340 5050 440 5060
rect 340 5030 370 5050
rect 410 5030 440 5050
rect 340 5020 440 5030
rect 510 5050 610 5060
rect 510 5030 540 5050
rect 580 5030 610 5050
rect 510 5020 610 5030
rect 680 5050 780 5060
rect 680 5030 710 5050
rect 750 5030 780 5050
rect 680 5020 780 5030
rect 850 5050 950 5060
rect 850 5030 880 5050
rect 920 5030 950 5050
rect 850 5020 950 5030
rect 1020 5050 1120 5060
rect 1020 5030 1050 5050
rect 1090 5030 1120 5050
rect 1020 5020 1120 5030
rect 1190 5050 1290 5060
rect 1190 5030 1220 5050
rect 1260 5030 1290 5050
rect 1190 5020 1290 5030
rect 1360 5050 1460 5060
rect 1360 5030 1390 5050
rect 1430 5030 1460 5050
rect 1360 5020 1460 5030
rect 1530 5050 1630 5060
rect 1530 5030 1560 5050
rect 1600 5030 1630 5050
rect 1530 5020 1630 5030
rect 1750 5050 1850 5060
rect 1750 5030 1780 5050
rect 1820 5030 1850 5050
rect 1750 5020 1850 5030
rect 1920 5050 2020 5060
rect 1920 5030 1950 5050
rect 1990 5030 2020 5050
rect 1920 5020 2020 5030
rect 2090 5050 2190 5060
rect 2090 5030 2120 5050
rect 2160 5030 2190 5050
rect 2090 5020 2190 5030
rect 2260 5050 2360 5060
rect 2260 5030 2290 5050
rect 2330 5030 2360 5050
rect 2260 5020 2360 5030
rect 2430 5050 2530 5060
rect 2430 5030 2460 5050
rect 2500 5030 2530 5050
rect 2430 5020 2530 5030
rect 2600 5050 2700 5060
rect 2600 5030 2630 5050
rect 2670 5030 2700 5050
rect 2600 5020 2700 5030
rect 2770 5050 2870 5060
rect 2770 5030 2800 5050
rect 2840 5030 2870 5050
rect 2770 5020 2870 5030
rect 2940 5050 3040 5060
rect 2940 5030 2970 5050
rect 3010 5030 3040 5050
rect 2940 5020 3040 5030
rect 3110 5050 3210 5060
rect 3110 5030 3140 5050
rect 3180 5030 3210 5050
rect 3110 5020 3210 5030
rect 3280 5050 3380 5060
rect 3280 5030 3310 5050
rect 3350 5030 3380 5050
rect 3280 5020 3380 5030
rect -280 4010 -80 4020
rect 0 4010 100 4020
rect 170 4010 270 4020
rect 340 4010 440 4020
rect 510 4010 610 4020
rect 680 4010 780 4020
rect 850 4010 950 4020
rect 1020 4010 1120 4020
rect 1190 4010 1290 4020
rect 1360 4010 1460 4020
rect 1530 4010 1630 4020
rect 1750 4010 1850 4020
rect 1920 4010 2020 4020
rect 2090 4010 2190 4020
rect 2260 4010 2360 4020
rect 2430 4010 2530 4020
rect 2600 4010 2700 4020
rect 2770 4010 2870 4020
rect 2940 4010 3040 4020
rect 3110 4010 3210 4020
rect 3280 4010 3380 4020
rect 3460 4010 3660 4020
rect -280 3990 -200 4010
rect -160 3990 30 4010
rect 70 3990 200 4010
rect 240 3990 370 4010
rect 410 3990 540 4010
rect 580 3990 710 4010
rect 750 3990 880 4010
rect 920 3990 1050 4010
rect 1090 3990 1220 4010
rect 1260 3990 1390 4010
rect 1430 3990 1560 4010
rect 1600 3990 1780 4010
rect 1820 3990 1950 4010
rect 1990 3990 2120 4010
rect 2160 3990 2290 4010
rect 2330 3990 2460 4010
rect 2500 3990 2630 4010
rect 2670 3990 2800 4010
rect 2840 3990 2970 4010
rect 3010 3990 3140 4010
rect 3180 3990 3310 4010
rect 3350 3990 3540 4010
rect 3580 3990 3660 4010
rect -280 3980 -80 3990
rect 0 3980 100 3990
rect 170 3980 270 3990
rect 340 3980 440 3990
rect 510 3980 610 3990
rect 680 3980 780 3990
rect 850 3980 950 3990
rect 1020 3980 1120 3990
rect 1190 3980 1290 3990
rect 1360 3980 1460 3990
rect 1530 3980 1630 3990
rect 1750 3980 1850 3990
rect 1920 3980 2020 3990
rect 2090 3980 2190 3990
rect 2260 3980 2360 3990
rect 2430 3980 2530 3990
rect 2600 3980 2700 3990
rect 2770 3980 2870 3990
rect 2940 3980 3040 3990
rect 3110 3980 3210 3990
rect 3280 3980 3380 3990
rect 3460 3980 3660 3990
rect -280 3470 -80 3480
rect -280 3450 -200 3470
rect -160 3450 -80 3470
rect -280 3440 -80 3450
rect 0 2970 100 2980
rect -280 2930 -80 2940
rect -280 2910 -200 2930
rect -160 2910 -80 2930
rect -280 2900 -80 2910
rect 0 2950 30 2970
rect 70 2950 100 2970
rect 0 2940 100 2950
rect 0 2870 100 2900
rect 170 2970 270 2980
rect 170 2950 200 2970
rect 240 2950 270 2970
rect 170 2940 270 2950
rect 170 2870 270 2900
rect 340 2970 440 2980
rect 340 2950 370 2970
rect 410 2950 440 2970
rect 340 2940 440 2950
rect 340 2870 440 2900
rect 510 2970 610 2980
rect 510 2950 540 2970
rect 580 2950 610 2970
rect 510 2940 610 2950
rect 510 2870 610 2900
rect 680 2970 780 2980
rect 680 2950 710 2970
rect 750 2950 780 2970
rect 680 2940 780 2950
rect 680 2870 780 2900
rect 850 2970 950 2980
rect 850 2950 880 2970
rect 920 2950 950 2970
rect 850 2940 950 2950
rect 850 2870 950 2900
rect 1020 2970 1120 2980
rect 1020 2950 1050 2970
rect 1090 2950 1120 2970
rect 1020 2940 1120 2950
rect 1020 2870 1120 2900
rect 1190 2970 1290 2980
rect 1190 2950 1220 2970
rect 1260 2950 1290 2970
rect 1190 2940 1290 2950
rect 1190 2870 1290 2900
rect 1360 2970 1460 2980
rect 1360 2950 1390 2970
rect 1430 2950 1460 2970
rect 1360 2940 1460 2950
rect 1360 2870 1460 2900
rect 1530 2970 1630 2980
rect 1530 2950 1560 2970
rect 1600 2950 1630 2970
rect 1530 2940 1630 2950
rect 1530 2870 1630 2900
rect 3460 3470 3660 3480
rect 3460 3450 3540 3470
rect 3580 3450 3660 3470
rect 3460 3440 3660 3450
rect 1750 2970 1850 2980
rect 1750 2950 1780 2970
rect 1820 2950 1850 2970
rect 1750 2940 1850 2950
rect 1750 2870 1850 2900
rect 1920 2970 2020 2980
rect 1920 2950 1950 2970
rect 1990 2950 2020 2970
rect 1920 2940 2020 2950
rect 1920 2870 2020 2900
rect 2090 2970 2190 2980
rect 2090 2950 2120 2970
rect 2160 2950 2190 2970
rect 2090 2940 2190 2950
rect 2090 2870 2190 2900
rect 2260 2970 2360 2980
rect 2260 2950 2290 2970
rect 2330 2950 2360 2970
rect 2260 2940 2360 2950
rect 2260 2870 2360 2900
rect 2430 2970 2530 2980
rect 2430 2950 2460 2970
rect 2500 2950 2530 2970
rect 2430 2940 2530 2950
rect 2430 2870 2530 2900
rect 2600 2970 2700 2980
rect 2600 2950 2630 2970
rect 2670 2950 2700 2970
rect 2600 2940 2700 2950
rect 2600 2870 2700 2900
rect 2770 2970 2870 2980
rect 2770 2950 2800 2970
rect 2840 2950 2870 2970
rect 2770 2940 2870 2950
rect 2770 2870 2870 2900
rect 2940 2970 3040 2980
rect 2940 2950 2970 2970
rect 3010 2950 3040 2970
rect 2940 2940 3040 2950
rect 2940 2870 3040 2900
rect 3110 2970 3210 2980
rect 3110 2950 3140 2970
rect 3180 2950 3210 2970
rect 3110 2940 3210 2950
rect 3110 2870 3210 2900
rect 3280 2970 3380 2980
rect 3280 2950 3310 2970
rect 3350 2950 3380 2970
rect 3280 2940 3380 2950
rect 3280 2870 3380 2900
rect 3460 2930 3660 2940
rect 3460 2910 3540 2930
rect 3580 2910 3660 2930
rect 3460 2900 3660 2910
rect 0 2760 100 2770
rect 0 2740 30 2760
rect 70 2740 100 2760
rect 0 2730 100 2740
rect 170 2760 270 2770
rect 170 2740 200 2760
rect 240 2740 270 2760
rect 170 2730 270 2740
rect 340 2760 440 2770
rect 340 2740 370 2760
rect 410 2740 440 2760
rect 340 2730 440 2740
rect 510 2760 610 2770
rect 510 2740 540 2760
rect 580 2740 610 2760
rect 510 2730 610 2740
rect 680 2760 780 2770
rect 680 2740 710 2760
rect 750 2740 780 2760
rect 680 2730 780 2740
rect 850 2760 950 2770
rect 850 2740 880 2760
rect 920 2740 950 2760
rect 850 2730 950 2740
rect 1020 2760 1120 2770
rect 1020 2740 1050 2760
rect 1090 2740 1120 2760
rect 1020 2730 1120 2740
rect 1190 2760 1290 2770
rect 1190 2740 1220 2760
rect 1260 2740 1290 2760
rect 1190 2730 1290 2740
rect 1360 2760 1460 2770
rect 1360 2740 1390 2760
rect 1430 2740 1460 2760
rect 1360 2730 1460 2740
rect 1530 2760 1630 2770
rect 1530 2740 1560 2760
rect 1600 2740 1630 2760
rect 1530 2730 1630 2740
rect 1750 2760 1850 2770
rect 1750 2740 1780 2760
rect 1820 2740 1850 2760
rect 1750 2730 1850 2740
rect 1920 2760 2020 2770
rect 1920 2740 1950 2760
rect 1990 2740 2020 2760
rect 1920 2730 2020 2740
rect 2090 2760 2190 2770
rect 2090 2740 2120 2760
rect 2160 2740 2190 2760
rect 2090 2730 2190 2740
rect 2260 2760 2360 2770
rect 2260 2740 2290 2760
rect 2330 2740 2360 2760
rect 2260 2730 2360 2740
rect 2430 2760 2530 2770
rect 2430 2740 2460 2760
rect 2500 2740 2530 2760
rect 2430 2730 2530 2740
rect 2600 2760 2700 2770
rect 2600 2740 2630 2760
rect 2670 2740 2700 2760
rect 2600 2730 2700 2740
rect 2770 2760 2870 2770
rect 2770 2740 2800 2760
rect 2840 2740 2870 2760
rect 2770 2730 2870 2740
rect 2940 2760 3040 2770
rect 2940 2740 2970 2760
rect 3010 2740 3040 2760
rect 2940 2730 3040 2740
rect 3110 2760 3210 2770
rect 3110 2740 3140 2760
rect 3180 2740 3210 2760
rect 3110 2730 3210 2740
rect 3280 2760 3380 2770
rect 3280 2740 3310 2760
rect 3350 2740 3380 2760
rect 3280 2730 3380 2740
rect 0 2280 100 2290
rect 0 2260 30 2280
rect 70 2260 100 2280
rect 0 2250 100 2260
rect 170 2280 270 2290
rect 170 2260 200 2280
rect 240 2260 270 2280
rect 170 2250 270 2260
rect 340 2280 440 2290
rect 340 2260 370 2280
rect 410 2260 440 2280
rect 340 2250 440 2260
rect 510 2280 610 2290
rect 510 2260 540 2280
rect 580 2260 610 2280
rect 510 2250 610 2260
rect 680 2280 780 2290
rect 680 2260 710 2280
rect 750 2260 780 2280
rect 680 2250 780 2260
rect 850 2280 950 2290
rect 850 2260 880 2280
rect 920 2260 950 2280
rect 850 2250 950 2260
rect 1020 2280 1120 2290
rect 1020 2260 1050 2280
rect 1090 2260 1120 2280
rect 1020 2250 1120 2260
rect 1190 2280 1290 2290
rect 1190 2260 1220 2280
rect 1260 2260 1290 2280
rect 1190 2250 1290 2260
rect 1360 2280 1460 2290
rect 1360 2260 1390 2280
rect 1430 2260 1460 2280
rect 1360 2250 1460 2260
rect 1530 2280 1630 2290
rect 1530 2260 1560 2280
rect 1600 2260 1630 2280
rect 1530 2250 1630 2260
rect 1750 2280 1850 2290
rect 1750 2260 1780 2280
rect 1820 2260 1850 2280
rect 1750 2250 1850 2260
rect 1920 2280 2020 2290
rect 1920 2260 1950 2280
rect 1990 2260 2020 2280
rect 1920 2250 2020 2260
rect 2090 2280 2190 2290
rect 2090 2260 2120 2280
rect 2160 2260 2190 2280
rect 2090 2250 2190 2260
rect 2260 2280 2360 2290
rect 2260 2260 2290 2280
rect 2330 2260 2360 2280
rect 2260 2250 2360 2260
rect 2430 2280 2530 2290
rect 2430 2260 2460 2280
rect 2500 2260 2530 2280
rect 2430 2250 2530 2260
rect 2600 2280 2700 2290
rect 2600 2260 2630 2280
rect 2670 2260 2700 2280
rect 2600 2250 2700 2260
rect 2770 2280 2870 2290
rect 2770 2260 2800 2280
rect 2840 2260 2870 2280
rect 2770 2250 2870 2260
rect 2940 2280 3040 2290
rect 2940 2260 2970 2280
rect 3010 2260 3040 2280
rect 2940 2250 3040 2260
rect 3110 2280 3210 2290
rect 3110 2260 3140 2280
rect 3180 2260 3210 2280
rect 3110 2250 3210 2260
rect 3280 2280 3380 2290
rect 3280 2260 3310 2280
rect 3350 2260 3380 2280
rect 3280 2250 3380 2260
rect -280 2110 -80 2120
rect -280 2090 -200 2110
rect -160 2090 -80 2110
rect -280 2080 -80 2090
rect 0 2120 100 2150
rect 0 2070 100 2080
rect 0 2050 30 2070
rect 70 2050 100 2070
rect 0 2040 100 2050
rect 170 2120 270 2150
rect 170 2070 270 2080
rect 170 2050 200 2070
rect 240 2050 270 2070
rect 170 2040 270 2050
rect 340 2120 440 2150
rect 340 2070 440 2080
rect 340 2050 370 2070
rect 410 2050 440 2070
rect 340 2040 440 2050
rect 510 2120 610 2150
rect 510 2070 610 2080
rect 510 2050 540 2070
rect 580 2050 610 2070
rect 510 2040 610 2050
rect 680 2120 780 2150
rect 680 2070 780 2080
rect 680 2050 710 2070
rect 750 2050 780 2070
rect 680 2040 780 2050
rect 850 2120 950 2150
rect 850 2070 950 2080
rect 850 2050 880 2070
rect 920 2050 950 2070
rect 850 2040 950 2050
rect 1020 2120 1120 2150
rect 1020 2070 1120 2080
rect 1020 2050 1050 2070
rect 1090 2050 1120 2070
rect 1020 2040 1120 2050
rect 1190 2120 1290 2150
rect 1190 2070 1290 2080
rect 1190 2050 1220 2070
rect 1260 2050 1290 2070
rect 1190 2040 1290 2050
rect 1360 2120 1460 2150
rect 1360 2070 1460 2080
rect 1360 2050 1390 2070
rect 1430 2050 1460 2070
rect 1360 2040 1460 2050
rect 1530 2120 1630 2150
rect 1530 2070 1630 2080
rect 1530 2050 1560 2070
rect 1600 2050 1630 2070
rect 1530 2040 1630 2050
rect -280 1570 -80 1580
rect -280 1550 -200 1570
rect -160 1550 -80 1570
rect -280 1540 -80 1550
rect 1750 2120 1850 2150
rect 1750 2070 1850 2080
rect 1750 2050 1780 2070
rect 1820 2050 1850 2070
rect 1750 2040 1850 2050
rect 1920 2120 2020 2150
rect 1920 2070 2020 2080
rect 1920 2050 1950 2070
rect 1990 2050 2020 2070
rect 1920 2040 2020 2050
rect 2090 2120 2190 2150
rect 2090 2070 2190 2080
rect 2090 2050 2120 2070
rect 2160 2050 2190 2070
rect 2090 2040 2190 2050
rect 2260 2120 2360 2150
rect 2260 2070 2360 2080
rect 2260 2050 2290 2070
rect 2330 2050 2360 2070
rect 2260 2040 2360 2050
rect 2430 2120 2530 2150
rect 2430 2070 2530 2080
rect 2430 2050 2460 2070
rect 2500 2050 2530 2070
rect 2430 2040 2530 2050
rect 2600 2120 2700 2150
rect 2600 2070 2700 2080
rect 2600 2050 2630 2070
rect 2670 2050 2700 2070
rect 2600 2040 2700 2050
rect 2770 2120 2870 2150
rect 2770 2070 2870 2080
rect 2770 2050 2800 2070
rect 2840 2050 2870 2070
rect 2770 2040 2870 2050
rect 2940 2120 3040 2150
rect 2940 2070 3040 2080
rect 2940 2050 2970 2070
rect 3010 2050 3040 2070
rect 2940 2040 3040 2050
rect 3110 2120 3210 2150
rect 3110 2070 3210 2080
rect 3110 2050 3140 2070
rect 3180 2050 3210 2070
rect 3110 2040 3210 2050
rect 3280 2120 3380 2150
rect 3280 2070 3380 2080
rect 3280 2050 3310 2070
rect 3350 2050 3380 2070
rect 3460 2110 3660 2120
rect 3460 2090 3540 2110
rect 3580 2090 3660 2110
rect 3460 2080 3660 2090
rect 3280 2040 3380 2050
rect 3460 1570 3660 1580
rect 3460 1550 3540 1570
rect 3580 1550 3660 1570
rect 3460 1540 3660 1550
rect -280 1030 -80 1040
rect 0 1030 100 1040
rect 170 1030 270 1040
rect 340 1030 440 1040
rect 510 1030 610 1040
rect 680 1030 780 1040
rect 850 1030 950 1040
rect 1020 1030 1120 1040
rect 1190 1030 1290 1040
rect 1360 1030 1460 1040
rect 1530 1030 1630 1040
rect 1750 1030 1850 1040
rect 1920 1030 2020 1040
rect 2090 1030 2190 1040
rect 2260 1030 2360 1040
rect 2430 1030 2530 1040
rect 2600 1030 2700 1040
rect 2770 1030 2870 1040
rect 2940 1030 3040 1040
rect 3110 1030 3210 1040
rect 3280 1030 3380 1040
rect 3460 1030 3660 1040
rect -280 1010 -200 1030
rect -160 1010 30 1030
rect 70 1010 200 1030
rect 240 1010 370 1030
rect 410 1010 540 1030
rect 580 1010 710 1030
rect 750 1010 880 1030
rect 920 1010 1050 1030
rect 1090 1010 1220 1030
rect 1260 1010 1390 1030
rect 1430 1010 1560 1030
rect 1600 1010 1780 1030
rect 1820 1010 1950 1030
rect 1990 1010 2120 1030
rect 2160 1010 2290 1030
rect 2330 1010 2460 1030
rect 2500 1010 2630 1030
rect 2670 1010 2800 1030
rect 2840 1010 2970 1030
rect 3010 1010 3140 1030
rect 3180 1010 3310 1030
rect 3350 1010 3540 1030
rect 3580 1010 3660 1030
rect -280 1000 -80 1010
rect 0 1000 100 1010
rect 170 1000 270 1010
rect 340 1000 440 1010
rect 510 1000 610 1010
rect 680 1000 780 1010
rect 850 1000 950 1010
rect 1020 1000 1120 1010
rect 1190 1000 1290 1010
rect 1360 1000 1460 1010
rect 1530 1000 1630 1010
rect 1750 1000 1850 1010
rect 1920 1000 2020 1010
rect 2090 1000 2190 1010
rect 2260 1000 2360 1010
rect 2430 1000 2530 1010
rect 2600 1000 2700 1010
rect 2770 1000 2870 1010
rect 2940 1000 3040 1010
rect 3110 1000 3210 1010
rect 3280 1000 3380 1010
rect 3460 1000 3660 1010
rect 0 -10 100 0
rect 0 -30 30 -10
rect 70 -30 100 -10
rect 0 -40 100 -30
rect 170 -10 270 0
rect 170 -30 200 -10
rect 240 -30 270 -10
rect 170 -40 270 -30
rect 340 -10 440 0
rect 340 -30 370 -10
rect 410 -30 440 -10
rect 340 -40 440 -30
rect 510 -10 610 0
rect 510 -30 540 -10
rect 580 -30 610 -10
rect 510 -40 610 -30
rect 680 -10 780 0
rect 680 -30 710 -10
rect 750 -30 780 -10
rect 680 -40 780 -30
rect 850 -10 950 0
rect 850 -30 880 -10
rect 920 -30 950 -10
rect 850 -40 950 -30
rect 1020 -10 1120 0
rect 1020 -30 1050 -10
rect 1090 -30 1120 -10
rect 1020 -40 1120 -30
rect 1190 -10 1290 0
rect 1190 -30 1220 -10
rect 1260 -30 1290 -10
rect 1190 -40 1290 -30
rect 1360 -10 1460 0
rect 1360 -30 1390 -10
rect 1430 -30 1460 -10
rect 1360 -40 1460 -30
rect 1530 -10 1630 0
rect 1530 -30 1560 -10
rect 1600 -30 1630 -10
rect 1530 -40 1630 -30
rect 1750 -10 1850 0
rect 1750 -30 1780 -10
rect 1820 -30 1850 -10
rect 1750 -40 1850 -30
rect 1920 -10 2020 0
rect 1920 -30 1950 -10
rect 1990 -30 2020 -10
rect 1920 -40 2020 -30
rect 2090 -10 2190 0
rect 2090 -30 2120 -10
rect 2160 -30 2190 -10
rect 2090 -40 2190 -30
rect 2260 -10 2360 0
rect 2260 -30 2290 -10
rect 2330 -30 2360 -10
rect 2260 -40 2360 -30
rect 2430 -10 2530 0
rect 2430 -30 2460 -10
rect 2500 -30 2530 -10
rect 2430 -40 2530 -30
rect 2600 -10 2700 0
rect 2600 -30 2630 -10
rect 2670 -30 2700 -10
rect 2600 -40 2700 -30
rect 2770 -10 2870 0
rect 2770 -30 2800 -10
rect 2840 -30 2870 -10
rect 2770 -40 2870 -30
rect 2940 -10 3040 0
rect 2940 -30 2970 -10
rect 3010 -30 3040 -10
rect 2940 -40 3040 -30
rect 3110 -10 3210 0
rect 3110 -30 3140 -10
rect 3180 -30 3210 -10
rect 3110 -40 3210 -30
rect 3280 -10 3380 0
rect 3280 -30 3310 -10
rect 3350 -30 3380 -10
rect 3280 -40 3380 -30
<< ndiffc >>
rect -190 2590 -170 2630
rect -50 2590 -30 2630
rect 90 2590 110 2630
rect 230 2590 250 2630
rect 370 2590 390 2630
rect 510 2590 530 2630
rect 650 2590 670 2630
rect 790 2590 810 2630
rect 930 2590 950 2630
rect 1070 2590 1090 2630
rect 1210 2590 1230 2630
rect 1560 2640 1580 2660
rect 1800 2640 1820 2660
rect 1350 2590 1370 2630
rect 1560 2570 1580 2590
rect 1800 2570 1820 2590
rect 2010 2590 2030 2630
rect 2150 2590 2170 2630
rect 2290 2590 2310 2630
rect 2430 2590 2450 2630
rect 2570 2590 2590 2630
rect 2710 2590 2730 2630
rect 2850 2590 2870 2630
rect 2990 2590 3010 2630
rect 3130 2590 3150 2630
rect 3270 2590 3290 2630
rect 3410 2590 3430 2630
rect 3550 2590 3570 2630
rect 1560 2500 1580 2520
rect 1800 2500 1820 2520
rect -190 2390 -170 2430
rect -50 2390 -30 2430
rect 90 2390 110 2430
rect 230 2390 250 2430
rect 370 2390 390 2430
rect 510 2390 530 2430
rect 650 2390 670 2430
rect 790 2390 810 2430
rect 930 2390 950 2430
rect 1070 2390 1090 2430
rect 1210 2390 1230 2430
rect 1350 2390 1370 2430
rect 1560 2430 1580 2450
rect 1800 2430 1820 2450
rect 2010 2390 2030 2430
rect 1560 2360 1580 2380
rect 1800 2360 1820 2380
rect 2150 2390 2170 2430
rect 2290 2390 2310 2430
rect 2430 2390 2450 2430
rect 2570 2390 2590 2430
rect 2710 2390 2730 2430
rect 2850 2390 2870 2430
rect 2990 2390 3010 2430
rect 3130 2390 3150 2430
rect 3270 2390 3290 2430
rect 3410 2390 3430 2430
rect 3550 2390 3570 2430
<< pdiffc >>
rect 30 5030 70 5050
rect 200 5030 240 5050
rect 370 5030 410 5050
rect 540 5030 580 5050
rect 710 5030 750 5050
rect 880 5030 920 5050
rect 1050 5030 1090 5050
rect 1220 5030 1260 5050
rect 1390 5030 1430 5050
rect 1560 5030 1600 5050
rect 1780 5030 1820 5050
rect 1950 5030 1990 5050
rect 2120 5030 2160 5050
rect 2290 5030 2330 5050
rect 2460 5030 2500 5050
rect 2630 5030 2670 5050
rect 2800 5030 2840 5050
rect 2970 5030 3010 5050
rect 3140 5030 3180 5050
rect 3310 5030 3350 5050
rect -200 3990 -160 4010
rect 30 3990 70 4010
rect 200 3990 240 4010
rect 370 3990 410 4010
rect 540 3990 580 4010
rect 710 3990 750 4010
rect 880 3990 920 4010
rect 1050 3990 1090 4010
rect 1220 3990 1260 4010
rect 1390 3990 1430 4010
rect 1560 3990 1600 4010
rect 1780 3990 1820 4010
rect 1950 3990 1990 4010
rect 2120 3990 2160 4010
rect 2290 3990 2330 4010
rect 2460 3990 2500 4010
rect 2630 3990 2670 4010
rect 2800 3990 2840 4010
rect 2970 3990 3010 4010
rect 3140 3990 3180 4010
rect 3310 3990 3350 4010
rect 3540 3990 3580 4010
rect -200 3450 -160 3470
rect -200 2910 -160 2930
rect 30 2950 70 2970
rect 200 2950 240 2970
rect 370 2950 410 2970
rect 540 2950 580 2970
rect 710 2950 750 2970
rect 880 2950 920 2970
rect 1050 2950 1090 2970
rect 1220 2950 1260 2970
rect 1390 2950 1430 2970
rect 1560 2950 1600 2970
rect 3540 3450 3580 3470
rect 1780 2950 1820 2970
rect 1950 2950 1990 2970
rect 2120 2950 2160 2970
rect 2290 2950 2330 2970
rect 2460 2950 2500 2970
rect 2630 2950 2670 2970
rect 2800 2950 2840 2970
rect 2970 2950 3010 2970
rect 3140 2950 3180 2970
rect 3310 2950 3350 2970
rect 3540 2910 3580 2930
rect 30 2740 70 2760
rect 200 2740 240 2760
rect 370 2740 410 2760
rect 540 2740 580 2760
rect 710 2740 750 2760
rect 880 2740 920 2760
rect 1050 2740 1090 2760
rect 1220 2740 1260 2760
rect 1390 2740 1430 2760
rect 1560 2740 1600 2760
rect 1780 2740 1820 2760
rect 1950 2740 1990 2760
rect 2120 2740 2160 2760
rect 2290 2740 2330 2760
rect 2460 2740 2500 2760
rect 2630 2740 2670 2760
rect 2800 2740 2840 2760
rect 2970 2740 3010 2760
rect 3140 2740 3180 2760
rect 3310 2740 3350 2760
rect 30 2260 70 2280
rect 200 2260 240 2280
rect 370 2260 410 2280
rect 540 2260 580 2280
rect 710 2260 750 2280
rect 880 2260 920 2280
rect 1050 2260 1090 2280
rect 1220 2260 1260 2280
rect 1390 2260 1430 2280
rect 1560 2260 1600 2280
rect 1780 2260 1820 2280
rect 1950 2260 1990 2280
rect 2120 2260 2160 2280
rect 2290 2260 2330 2280
rect 2460 2260 2500 2280
rect 2630 2260 2670 2280
rect 2800 2260 2840 2280
rect 2970 2260 3010 2280
rect 3140 2260 3180 2280
rect 3310 2260 3350 2280
rect -200 2090 -160 2110
rect 30 2050 70 2070
rect 200 2050 240 2070
rect 370 2050 410 2070
rect 540 2050 580 2070
rect 710 2050 750 2070
rect 880 2050 920 2070
rect 1050 2050 1090 2070
rect 1220 2050 1260 2070
rect 1390 2050 1430 2070
rect 1560 2050 1600 2070
rect -200 1550 -160 1570
rect 1780 2050 1820 2070
rect 1950 2050 1990 2070
rect 2120 2050 2160 2070
rect 2290 2050 2330 2070
rect 2460 2050 2500 2070
rect 2630 2050 2670 2070
rect 2800 2050 2840 2070
rect 2970 2050 3010 2070
rect 3140 2050 3180 2070
rect 3310 2050 3350 2070
rect 3540 2090 3580 2110
rect 3540 1550 3580 1570
rect -200 1010 -160 1030
rect 30 1010 70 1030
rect 200 1010 240 1030
rect 370 1010 410 1030
rect 540 1010 580 1030
rect 710 1010 750 1030
rect 880 1010 920 1030
rect 1050 1010 1090 1030
rect 1220 1010 1260 1030
rect 1390 1010 1430 1030
rect 1560 1010 1600 1030
rect 1780 1010 1820 1030
rect 1950 1010 1990 1030
rect 2120 1010 2160 1030
rect 2290 1010 2330 1030
rect 2460 1010 2500 1030
rect 2630 1010 2670 1030
rect 2800 1010 2840 1030
rect 2970 1010 3010 1030
rect 3140 1010 3180 1030
rect 3310 1010 3350 1030
rect 3540 1010 3580 1030
rect 30 -30 70 -10
rect 200 -30 240 -10
rect 370 -30 410 -10
rect 540 -30 580 -10
rect 710 -30 750 -10
rect 880 -30 920 -10
rect 1050 -30 1090 -10
rect 1220 -30 1260 -10
rect 1390 -30 1430 -10
rect 1560 -30 1600 -10
rect 1780 -30 1820 -10
rect 1950 -30 1990 -10
rect 2120 -30 2160 -10
rect 2290 -30 2330 -10
rect 2460 -30 2500 -10
rect 2630 -30 2670 -10
rect 2800 -30 2840 -10
rect 2970 -30 3010 -10
rect 3140 -30 3180 -10
rect 3310 -30 3350 -10
<< psubdiff >>
rect -240 2630 -200 2650
rect -240 2590 -230 2630
rect -210 2590 -200 2630
rect -240 2560 -200 2590
rect 3580 2630 3620 2650
rect 3580 2590 3590 2630
rect 3610 2590 3620 2630
rect 3580 2560 3620 2590
rect 1400 2520 1460 2540
rect 1400 2500 1420 2520
rect 1440 2500 1460 2520
rect 1400 2480 1460 2500
rect 1920 2520 1980 2540
rect 1920 2500 1940 2520
rect 1960 2500 1980 2520
rect 1920 2480 1980 2500
rect -240 2430 -200 2460
rect -240 2390 -230 2430
rect -210 2390 -200 2430
rect -240 2370 -200 2390
rect 3580 2430 3620 2460
rect 3580 2390 3590 2430
rect 3610 2390 3620 2430
rect 3580 2370 3620 2390
<< nsubdiff >>
rect 0 5070 30 5090
rect 70 5070 100 5090
rect 0 5060 100 5070
rect 170 5070 200 5090
rect 240 5070 270 5090
rect 170 5060 270 5070
rect 340 5070 370 5090
rect 410 5070 440 5090
rect 340 5060 440 5070
rect 510 5070 540 5090
rect 580 5070 610 5090
rect 510 5060 610 5070
rect 680 5070 710 5090
rect 750 5070 780 5090
rect 680 5060 780 5070
rect 850 5070 880 5090
rect 920 5070 950 5090
rect 850 5060 950 5070
rect 1020 5070 1050 5090
rect 1090 5070 1120 5090
rect 1020 5060 1120 5070
rect 1190 5070 1220 5090
rect 1260 5070 1290 5090
rect 1190 5060 1290 5070
rect 1360 5070 1390 5090
rect 1430 5070 1460 5090
rect 1360 5060 1460 5070
rect 1530 5070 1560 5090
rect 1600 5070 1630 5090
rect 1530 5060 1630 5070
rect 1750 5070 1780 5090
rect 1820 5070 1850 5090
rect 1750 5060 1850 5070
rect 1920 5070 1950 5090
rect 1990 5070 2020 5090
rect 1920 5060 2020 5070
rect 2090 5070 2120 5090
rect 2160 5070 2190 5090
rect 2090 5060 2190 5070
rect 2260 5070 2290 5090
rect 2330 5070 2360 5090
rect 2260 5060 2360 5070
rect 2430 5070 2460 5090
rect 2500 5070 2530 5090
rect 2430 5060 2530 5070
rect 2600 5070 2630 5090
rect 2670 5070 2700 5090
rect 2600 5060 2700 5070
rect 2770 5070 2800 5090
rect 2840 5070 2870 5090
rect 2770 5060 2870 5070
rect 2940 5070 2970 5090
rect 3010 5070 3040 5090
rect 2940 5060 3040 5070
rect 3110 5070 3140 5090
rect 3180 5070 3210 5090
rect 3110 5060 3210 5070
rect 3280 5070 3310 5090
rect 3350 5070 3380 5090
rect 3280 5060 3380 5070
rect 0 2930 100 2940
rect 0 2910 30 2930
rect 70 2910 100 2930
rect 0 2900 100 2910
rect 170 2930 270 2940
rect 170 2910 200 2930
rect 240 2910 270 2930
rect 170 2900 270 2910
rect 340 2930 440 2940
rect 340 2910 370 2930
rect 410 2910 440 2930
rect 340 2900 440 2910
rect 510 2930 610 2940
rect 510 2910 540 2930
rect 580 2910 610 2930
rect 510 2900 610 2910
rect 680 2930 780 2940
rect 680 2910 710 2930
rect 750 2910 780 2930
rect 680 2900 780 2910
rect 850 2930 950 2940
rect 850 2910 880 2930
rect 920 2910 950 2930
rect 850 2900 950 2910
rect 1020 2930 1120 2940
rect 1020 2910 1050 2930
rect 1090 2910 1120 2930
rect 1020 2900 1120 2910
rect 1190 2930 1290 2940
rect 1190 2910 1220 2930
rect 1260 2910 1290 2930
rect 1190 2900 1290 2910
rect 1360 2930 1460 2940
rect 1360 2910 1390 2930
rect 1430 2910 1460 2930
rect 1360 2900 1460 2910
rect 1530 2930 1630 2940
rect 1530 2910 1560 2930
rect 1600 2910 1630 2930
rect 1530 2900 1630 2910
rect 1750 2930 1850 2940
rect 1750 2910 1780 2930
rect 1820 2910 1850 2930
rect 1750 2900 1850 2910
rect 1920 2930 2020 2940
rect 1920 2910 1950 2930
rect 1990 2910 2020 2930
rect 1920 2900 2020 2910
rect 2090 2930 2190 2940
rect 2090 2910 2120 2930
rect 2160 2910 2190 2930
rect 2090 2900 2190 2910
rect 2260 2930 2360 2940
rect 2260 2910 2290 2930
rect 2330 2910 2360 2930
rect 2260 2900 2360 2910
rect 2430 2930 2530 2940
rect 2430 2910 2460 2930
rect 2500 2910 2530 2930
rect 2430 2900 2530 2910
rect 2600 2930 2700 2940
rect 2600 2910 2630 2930
rect 2670 2910 2700 2930
rect 2600 2900 2700 2910
rect 2770 2930 2870 2940
rect 2770 2910 2800 2930
rect 2840 2910 2870 2930
rect 2770 2900 2870 2910
rect 2940 2930 3040 2940
rect 2940 2910 2970 2930
rect 3010 2910 3040 2930
rect 2940 2900 3040 2910
rect 3110 2930 3210 2940
rect 3110 2910 3140 2930
rect 3180 2910 3210 2930
rect 3110 2900 3210 2910
rect 3280 2930 3380 2940
rect 3280 2910 3310 2930
rect 3350 2910 3380 2930
rect 3280 2900 3380 2910
rect 0 2110 100 2120
rect 0 2090 30 2110
rect 70 2090 100 2110
rect 0 2080 100 2090
rect 170 2110 270 2120
rect 170 2090 200 2110
rect 240 2090 270 2110
rect 170 2080 270 2090
rect 340 2110 440 2120
rect 340 2090 370 2110
rect 410 2090 440 2110
rect 340 2080 440 2090
rect 510 2110 610 2120
rect 510 2090 540 2110
rect 580 2090 610 2110
rect 510 2080 610 2090
rect 680 2110 780 2120
rect 680 2090 710 2110
rect 750 2090 780 2110
rect 680 2080 780 2090
rect 850 2110 950 2120
rect 850 2090 880 2110
rect 920 2090 950 2110
rect 850 2080 950 2090
rect 1020 2110 1120 2120
rect 1020 2090 1050 2110
rect 1090 2090 1120 2110
rect 1020 2080 1120 2090
rect 1190 2110 1290 2120
rect 1190 2090 1220 2110
rect 1260 2090 1290 2110
rect 1190 2080 1290 2090
rect 1360 2110 1460 2120
rect 1360 2090 1390 2110
rect 1430 2090 1460 2110
rect 1360 2080 1460 2090
rect 1530 2110 1630 2120
rect 1530 2090 1560 2110
rect 1600 2090 1630 2110
rect 1530 2080 1630 2090
rect 1750 2110 1850 2120
rect 1750 2090 1780 2110
rect 1820 2090 1850 2110
rect 1750 2080 1850 2090
rect 1920 2110 2020 2120
rect 1920 2090 1950 2110
rect 1990 2090 2020 2110
rect 1920 2080 2020 2090
rect 2090 2110 2190 2120
rect 2090 2090 2120 2110
rect 2160 2090 2190 2110
rect 2090 2080 2190 2090
rect 2260 2110 2360 2120
rect 2260 2090 2290 2110
rect 2330 2090 2360 2110
rect 2260 2080 2360 2090
rect 2430 2110 2530 2120
rect 2430 2090 2460 2110
rect 2500 2090 2530 2110
rect 2430 2080 2530 2090
rect 2600 2110 2700 2120
rect 2600 2090 2630 2110
rect 2670 2090 2700 2110
rect 2600 2080 2700 2090
rect 2770 2110 2870 2120
rect 2770 2090 2800 2110
rect 2840 2090 2870 2110
rect 2770 2080 2870 2090
rect 2940 2110 3040 2120
rect 2940 2090 2970 2110
rect 3010 2090 3040 2110
rect 2940 2080 3040 2090
rect 3110 2110 3210 2120
rect 3110 2090 3140 2110
rect 3180 2090 3210 2110
rect 3110 2080 3210 2090
rect 3280 2110 3380 2120
rect 3280 2090 3310 2110
rect 3350 2090 3380 2110
rect 3280 2080 3380 2090
rect 0 -50 100 -40
rect 0 -70 30 -50
rect 70 -70 100 -50
rect 170 -50 270 -40
rect 170 -70 200 -50
rect 240 -70 270 -50
rect 340 -50 440 -40
rect 340 -70 370 -50
rect 410 -70 440 -50
rect 510 -50 610 -40
rect 510 -70 540 -50
rect 580 -70 610 -50
rect 680 -50 780 -40
rect 680 -70 710 -50
rect 750 -70 780 -50
rect 850 -50 950 -40
rect 850 -70 880 -50
rect 920 -70 950 -50
rect 1020 -50 1120 -40
rect 1020 -70 1050 -50
rect 1090 -70 1120 -50
rect 1190 -50 1290 -40
rect 1190 -70 1220 -50
rect 1260 -70 1290 -50
rect 1360 -50 1460 -40
rect 1360 -70 1390 -50
rect 1430 -70 1460 -50
rect 1530 -50 1630 -40
rect 1530 -70 1560 -50
rect 1600 -70 1630 -50
rect 1750 -50 1850 -40
rect 1750 -70 1780 -50
rect 1820 -70 1850 -50
rect 1920 -50 2020 -40
rect 1920 -70 1950 -50
rect 1990 -70 2020 -50
rect 2090 -50 2190 -40
rect 2090 -70 2120 -50
rect 2160 -70 2190 -50
rect 2260 -50 2360 -40
rect 2260 -70 2290 -50
rect 2330 -70 2360 -50
rect 2430 -50 2530 -40
rect 2430 -70 2460 -50
rect 2500 -70 2530 -50
rect 2600 -50 2700 -40
rect 2600 -70 2630 -50
rect 2670 -70 2700 -50
rect 2770 -50 2870 -40
rect 2770 -70 2800 -50
rect 2840 -70 2870 -50
rect 2940 -50 3040 -40
rect 2940 -70 2970 -50
rect 3010 -70 3040 -50
rect 3110 -50 3210 -40
rect 3110 -70 3140 -50
rect 3180 -70 3210 -50
rect 3280 -50 3380 -40
rect 3280 -70 3310 -50
rect 3350 -70 3380 -50
<< psubdiffcont >>
rect -230 2590 -210 2630
rect 3590 2590 3610 2630
rect 1420 2500 1440 2520
rect 1940 2500 1960 2520
rect -230 2390 -210 2430
rect 3590 2390 3610 2430
<< nsubdiffcont >>
rect 30 5070 70 5090
rect 200 5070 240 5090
rect 370 5070 410 5090
rect 540 5070 580 5090
rect 710 5070 750 5090
rect 880 5070 920 5090
rect 1050 5070 1090 5090
rect 1220 5070 1260 5090
rect 1390 5070 1430 5090
rect 1560 5070 1600 5090
rect 1780 5070 1820 5090
rect 1950 5070 1990 5090
rect 2120 5070 2160 5090
rect 2290 5070 2330 5090
rect 2460 5070 2500 5090
rect 2630 5070 2670 5090
rect 2800 5070 2840 5090
rect 2970 5070 3010 5090
rect 3140 5070 3180 5090
rect 3310 5070 3350 5090
rect 30 2910 70 2930
rect 200 2910 240 2930
rect 370 2910 410 2930
rect 540 2910 580 2930
rect 710 2910 750 2930
rect 880 2910 920 2930
rect 1050 2910 1090 2930
rect 1220 2910 1260 2930
rect 1390 2910 1430 2930
rect 1560 2910 1600 2930
rect 1780 2910 1820 2930
rect 1950 2910 1990 2930
rect 2120 2910 2160 2930
rect 2290 2910 2330 2930
rect 2460 2910 2500 2930
rect 2630 2910 2670 2930
rect 2800 2910 2840 2930
rect 2970 2910 3010 2930
rect 3140 2910 3180 2930
rect 3310 2910 3350 2930
rect 30 2090 70 2110
rect 200 2090 240 2110
rect 370 2090 410 2110
rect 540 2090 580 2110
rect 710 2090 750 2110
rect 880 2090 920 2110
rect 1050 2090 1090 2110
rect 1220 2090 1260 2110
rect 1390 2090 1430 2110
rect 1560 2090 1600 2110
rect 1780 2090 1820 2110
rect 1950 2090 1990 2110
rect 2120 2090 2160 2110
rect 2290 2090 2330 2110
rect 2460 2090 2500 2110
rect 2630 2090 2670 2110
rect 2800 2090 2840 2110
rect 2970 2090 3010 2110
rect 3140 2090 3180 2110
rect 3310 2090 3350 2110
rect 30 -70 70 -50
rect 200 -70 240 -50
rect 370 -70 410 -50
rect 540 -70 580 -50
rect 710 -70 750 -50
rect 880 -70 920 -50
rect 1050 -70 1090 -50
rect 1220 -70 1260 -50
rect 1390 -70 1430 -50
rect 1560 -70 1600 -50
rect 1780 -70 1820 -50
rect 1950 -70 1990 -50
rect 2120 -70 2160 -50
rect 2290 -70 2330 -50
rect 2460 -70 2500 -50
rect 2630 -70 2670 -50
rect 2800 -70 2840 -50
rect 2970 -70 3010 -50
rect 3140 -70 3180 -50
rect 3310 -70 3350 -50
<< poly >>
rect -60 5070 -20 5080
rect -60 5050 -50 5070
rect -30 5050 -20 5070
rect -60 5040 -20 5050
rect -40 5020 -20 5040
rect 3400 5070 3440 5080
rect 3400 5050 3410 5070
rect 3430 5050 3440 5070
rect 3400 5040 3440 5050
rect 3400 5020 3420 5040
rect -40 5000 0 5020
rect -310 4070 -270 4080
rect -310 4050 -300 4070
rect -280 4050 -270 4070
rect -310 4040 -270 4050
rect -310 3980 -290 4040
rect -20 4020 0 5000
rect 100 4530 120 5020
rect 150 4530 170 5020
rect 100 4510 170 4530
rect 100 4020 120 4510
rect 150 4020 170 4510
rect 270 4530 290 5020
rect 320 4530 340 5020
rect 270 4510 340 4530
rect 270 4020 290 4510
rect 320 4020 340 4510
rect 440 4530 460 5020
rect 490 4530 510 5020
rect 440 4510 510 4530
rect 440 4020 460 4510
rect 490 4020 510 4510
rect 610 4530 630 5020
rect 660 4530 680 5020
rect 610 4510 680 4530
rect 610 4020 630 4510
rect 660 4020 680 4510
rect 780 4530 800 5020
rect 830 4530 850 5020
rect 780 4510 850 4530
rect 780 4020 800 4510
rect 830 4020 850 4510
rect 950 4530 970 5020
rect 1000 4530 1020 5020
rect 950 4510 1020 4530
rect 950 4020 970 4510
rect 1000 4020 1020 4510
rect 1120 4530 1140 5020
rect 1170 4530 1190 5020
rect 1120 4510 1190 4530
rect 1120 4020 1140 4510
rect 1170 4020 1190 4510
rect 1290 4530 1310 5020
rect 1340 4530 1360 5020
rect 1290 4510 1360 4530
rect 1290 4020 1310 4510
rect 1340 4020 1360 4510
rect 1460 4530 1480 5020
rect 1510 4530 1530 5020
rect 1460 4510 1530 4530
rect 1460 4020 1480 4510
rect 1510 4020 1530 4510
rect 1630 4530 1650 5020
rect 1730 4530 1750 5020
rect 1630 4510 1750 4530
rect 1630 4020 1650 4510
rect 1730 4020 1750 4510
rect 1850 4530 1870 5020
rect 1900 4530 1920 5020
rect 1850 4510 1920 4530
rect 1850 4020 1870 4510
rect 1900 4020 1920 4510
rect 2020 4530 2040 5020
rect 2070 4530 2090 5020
rect 2020 4510 2090 4530
rect 2020 4020 2040 4510
rect 2070 4020 2090 4510
rect 2190 4530 2210 5020
rect 2240 4530 2260 5020
rect 2190 4510 2260 4530
rect 2190 4020 2210 4510
rect 2240 4020 2260 4510
rect 2360 4530 2380 5020
rect 2410 4530 2430 5020
rect 2360 4510 2430 4530
rect 2360 4020 2380 4510
rect 2410 4020 2430 4510
rect 2530 4530 2550 5020
rect 2580 4530 2600 5020
rect 2530 4510 2600 4530
rect 2530 4020 2550 4510
rect 2580 4020 2600 4510
rect 2700 4530 2720 5020
rect 2750 4530 2770 5020
rect 2700 4510 2770 4530
rect 2700 4020 2720 4510
rect 2750 4020 2770 4510
rect 2870 4530 2890 5020
rect 2920 4530 2940 5020
rect 2870 4510 2940 4530
rect 2870 4020 2890 4510
rect 2920 4020 2940 4510
rect 3040 4530 3060 5020
rect 3090 4530 3110 5020
rect 3040 4510 3110 4530
rect 3040 4020 3060 4510
rect 3090 4020 3110 4510
rect 3210 4530 3230 5020
rect 3260 4530 3280 5020
rect 3210 4510 3280 4530
rect 3210 4020 3230 4510
rect 3260 4020 3280 4510
rect 3380 5000 3420 5020
rect 3380 4020 3400 5000
rect 3650 4070 3690 4080
rect 3650 4050 3660 4070
rect 3680 4050 3690 4070
rect 3650 4040 3690 4050
rect 3670 3980 3690 4040
rect -310 3960 -280 3980
rect -300 3480 -280 3960
rect -80 3480 -60 3980
rect -300 2940 -280 3440
rect -80 2960 -60 3440
rect -20 2980 0 3980
rect 100 3490 120 3980
rect 150 3490 170 3980
rect 100 3470 170 3490
rect 100 2980 120 3470
rect 150 2980 170 3470
rect 270 3490 290 3980
rect 320 3490 340 3980
rect 270 3470 340 3490
rect 270 2980 290 3470
rect 320 2980 340 3470
rect 440 3490 460 3980
rect 490 3490 510 3980
rect 440 3470 510 3490
rect 440 2980 460 3470
rect 490 2980 510 3470
rect 610 3490 630 3980
rect 660 3490 680 3980
rect 610 3470 680 3490
rect 610 2980 630 3470
rect 660 2980 680 3470
rect 780 3490 800 3980
rect 830 3490 850 3980
rect 780 3470 850 3490
rect 780 2980 800 3470
rect 830 2980 850 3470
rect 950 3490 970 3980
rect 1000 3490 1020 3980
rect 950 3470 1020 3490
rect 950 2980 970 3470
rect 1000 2980 1020 3470
rect 1120 3490 1140 3980
rect 1170 3490 1190 3980
rect 1120 3470 1190 3490
rect 1120 2980 1140 3470
rect 1170 2980 1190 3470
rect 1290 3490 1310 3980
rect 1340 3490 1360 3980
rect 1290 3470 1360 3490
rect 1290 2980 1310 3470
rect 1340 2980 1360 3470
rect 1460 3490 1480 3980
rect 1510 3490 1530 3980
rect 1460 3470 1530 3490
rect 1460 2980 1480 3470
rect 1510 2980 1530 3470
rect 1630 3490 1650 3980
rect 1730 3490 1750 3980
rect 1630 3470 1750 3490
rect 1630 2980 1650 3470
rect -80 2940 -50 2960
rect -70 2880 -50 2940
rect -90 2870 -50 2880
rect -90 2850 -80 2870
rect -60 2850 -50 2870
rect -90 2840 -50 2850
rect -20 2770 0 2870
rect 100 2830 120 2870
rect 150 2830 170 2870
rect 100 2810 170 2830
rect 100 2770 120 2810
rect 150 2770 170 2810
rect 270 2830 290 2870
rect 320 2830 340 2870
rect 270 2810 340 2830
rect 270 2770 290 2810
rect 320 2770 340 2810
rect 440 2830 460 2870
rect 490 2830 510 2870
rect 440 2810 510 2830
rect 440 2770 460 2810
rect 490 2770 510 2810
rect 610 2830 630 2870
rect 660 2830 680 2870
rect 610 2810 680 2830
rect 610 2770 630 2810
rect 660 2770 680 2810
rect 780 2830 800 2870
rect 830 2830 850 2870
rect 780 2810 850 2830
rect 780 2770 800 2810
rect 830 2770 850 2810
rect 950 2830 970 2870
rect 1000 2830 1020 2870
rect 950 2810 1020 2830
rect 950 2770 970 2810
rect 1000 2770 1020 2810
rect 1120 2830 1140 2870
rect 1170 2830 1190 2870
rect 1120 2810 1190 2830
rect 1120 2770 1140 2810
rect 1170 2770 1190 2810
rect 1290 2830 1310 2870
rect 1340 2830 1360 2870
rect 1290 2810 1360 2830
rect 1290 2770 1310 2810
rect 1340 2770 1360 2810
rect 1460 2830 1480 2870
rect 1510 2830 1530 2870
rect 1460 2810 1530 2830
rect 1460 2770 1480 2810
rect 1510 2770 1530 2810
rect 1630 2830 1650 2870
rect 1680 2830 1700 3470
rect 1730 2980 1750 3470
rect 1850 3490 1870 3980
rect 1900 3490 1920 3980
rect 1850 3470 1920 3490
rect 1850 2980 1870 3470
rect 1900 2980 1920 3470
rect 2020 3490 2040 3980
rect 2070 3490 2090 3980
rect 2020 3470 2090 3490
rect 2020 2980 2040 3470
rect 2070 2980 2090 3470
rect 2190 3490 2210 3980
rect 2240 3490 2260 3980
rect 2190 3470 2260 3490
rect 2190 2980 2210 3470
rect 2240 2980 2260 3470
rect 2360 3490 2380 3980
rect 2410 3490 2430 3980
rect 2360 3470 2430 3490
rect 2360 2980 2380 3470
rect 2410 2980 2430 3470
rect 2530 3490 2550 3980
rect 2580 3490 2600 3980
rect 2530 3470 2600 3490
rect 2530 2980 2550 3470
rect 2580 2980 2600 3470
rect 2700 3490 2720 3980
rect 2750 3490 2770 3980
rect 2700 3470 2770 3490
rect 2700 2980 2720 3470
rect 2750 2980 2770 3470
rect 2870 3490 2890 3980
rect 2920 3490 2940 3980
rect 2870 3470 2940 3490
rect 2870 2980 2890 3470
rect 2920 2980 2940 3470
rect 3040 3490 3060 3980
rect 3090 3490 3110 3980
rect 3040 3470 3110 3490
rect 3040 2980 3060 3470
rect 3090 2980 3110 3470
rect 3210 3490 3230 3980
rect 3260 3490 3280 3980
rect 3210 3470 3280 3490
rect 3210 2980 3230 3470
rect 3260 2980 3280 3470
rect 3380 2980 3400 3980
rect 3440 3480 3460 3980
rect 3660 3960 3690 3980
rect 3660 3480 3680 3960
rect 3440 2960 3460 3440
rect 3430 2940 3460 2960
rect 3660 2940 3680 3440
rect 3430 2880 3450 2940
rect 3430 2870 3470 2880
rect 1730 2830 1750 2870
rect 1630 2810 1750 2830
rect 1630 2770 1660 2810
rect 1640 2710 1660 2770
rect -200 2700 -160 2710
rect -200 2680 -190 2700
rect -170 2690 -160 2700
rect 80 2700 120 2710
rect 80 2690 90 2700
rect -170 2680 -140 2690
rect 60 2680 90 2690
rect 110 2690 120 2700
rect 360 2700 400 2710
rect 360 2690 370 2700
rect 110 2680 140 2690
rect 340 2680 370 2690
rect 390 2690 400 2700
rect 640 2700 680 2710
rect 640 2690 650 2700
rect 390 2680 420 2690
rect 620 2680 650 2690
rect 670 2690 680 2700
rect 920 2700 960 2710
rect 920 2690 930 2700
rect 670 2680 700 2690
rect 900 2680 930 2690
rect 950 2690 960 2700
rect 1200 2700 1240 2710
rect 1200 2690 1210 2700
rect 950 2680 980 2690
rect 1180 2680 1210 2690
rect 1230 2690 1240 2700
rect 1610 2700 1660 2710
rect 1230 2680 1260 2690
rect 1610 2680 1620 2700
rect 1640 2680 1660 2700
rect -200 2670 -60 2680
rect -160 2660 -60 2670
rect -20 2670 220 2680
rect -20 2660 80 2670
rect 120 2660 220 2670
rect 260 2670 500 2680
rect 260 2660 360 2670
rect 400 2660 500 2670
rect 540 2670 780 2680
rect 540 2660 640 2670
rect 680 2660 780 2670
rect 820 2670 1060 2680
rect 820 2660 920 2670
rect 960 2660 1060 2670
rect 1100 2670 1340 2680
rect 1610 2670 1660 2680
rect 1720 2770 1750 2810
rect 1850 2830 1870 2870
rect 1900 2830 1920 2870
rect 1850 2810 1920 2830
rect 1850 2770 1870 2810
rect 1900 2770 1920 2810
rect 2020 2830 2040 2870
rect 2070 2830 2090 2870
rect 2020 2810 2090 2830
rect 2020 2770 2040 2810
rect 2070 2770 2090 2810
rect 2190 2830 2210 2870
rect 2240 2830 2260 2870
rect 2190 2810 2260 2830
rect 2190 2770 2210 2810
rect 2240 2770 2260 2810
rect 2360 2830 2380 2870
rect 2410 2830 2430 2870
rect 2360 2810 2430 2830
rect 2360 2770 2380 2810
rect 2410 2770 2430 2810
rect 2530 2830 2550 2870
rect 2580 2830 2600 2870
rect 2530 2810 2600 2830
rect 2530 2770 2550 2810
rect 2580 2770 2600 2810
rect 2700 2830 2720 2870
rect 2750 2830 2770 2870
rect 2700 2810 2770 2830
rect 2700 2770 2720 2810
rect 2750 2770 2770 2810
rect 2870 2830 2890 2870
rect 2920 2830 2940 2870
rect 2870 2810 2940 2830
rect 2870 2770 2890 2810
rect 2920 2770 2940 2810
rect 3040 2830 3060 2870
rect 3090 2830 3110 2870
rect 3040 2810 3110 2830
rect 3040 2770 3060 2810
rect 3090 2770 3110 2810
rect 3210 2830 3230 2870
rect 3260 2830 3280 2870
rect 3210 2810 3280 2830
rect 3210 2770 3230 2810
rect 3260 2770 3280 2810
rect 3380 2770 3400 2870
rect 3430 2850 3440 2870
rect 3460 2850 3470 2870
rect 3430 2840 3470 2850
rect 1720 2710 1740 2770
rect 1720 2700 1770 2710
rect 1720 2680 1740 2700
rect 1760 2680 1770 2700
rect 2140 2700 2180 2710
rect 2140 2690 2150 2700
rect 2120 2680 2150 2690
rect 2170 2690 2180 2700
rect 2420 2700 2460 2710
rect 2420 2690 2430 2700
rect 2170 2680 2200 2690
rect 2400 2680 2430 2690
rect 2450 2690 2460 2700
rect 2700 2700 2740 2710
rect 2700 2690 2710 2700
rect 2450 2680 2480 2690
rect 2680 2680 2710 2690
rect 2730 2690 2740 2700
rect 2980 2700 3020 2710
rect 2980 2690 2990 2700
rect 2730 2680 2760 2690
rect 2960 2680 2990 2690
rect 3010 2690 3020 2700
rect 3260 2700 3300 2710
rect 3260 2690 3270 2700
rect 3010 2680 3040 2690
rect 3240 2680 3270 2690
rect 3290 2690 3300 2700
rect 3540 2700 3580 2710
rect 3540 2690 3550 2700
rect 3290 2680 3320 2690
rect 3520 2680 3550 2690
rect 3570 2680 3580 2700
rect 1720 2670 1770 2680
rect 2040 2670 2280 2680
rect 1100 2660 1200 2670
rect 1240 2660 1340 2670
rect 2040 2660 2140 2670
rect 2180 2660 2280 2670
rect 2320 2670 2560 2680
rect 2320 2660 2420 2670
rect 2460 2660 2560 2670
rect 2600 2670 2840 2680
rect 2600 2660 2700 2670
rect 2740 2660 2840 2670
rect 2880 2670 3120 2680
rect 2880 2660 2980 2670
rect 3020 2660 3120 2670
rect 3160 2670 3400 2680
rect 3160 2660 3260 2670
rect 3300 2660 3400 2670
rect 3440 2670 3580 2680
rect 3440 2660 3540 2670
rect -160 2540 -60 2560
rect -20 2540 80 2560
rect 120 2540 220 2560
rect 260 2540 360 2560
rect 400 2540 500 2560
rect 540 2540 640 2560
rect 680 2540 780 2560
rect 820 2540 920 2560
rect 960 2540 1060 2560
rect 1100 2540 1200 2560
rect -160 2460 -60 2480
rect -20 2460 80 2480
rect 120 2460 220 2480
rect 260 2460 360 2480
rect 400 2460 500 2480
rect 540 2460 640 2480
rect 680 2460 780 2480
rect 820 2460 920 2480
rect 960 2460 1060 2480
rect 1100 2460 1200 2480
rect 1240 2540 1340 2560
rect 1240 2460 1340 2480
rect 2040 2540 2140 2560
rect 2040 2460 2140 2480
rect 2180 2540 2280 2560
rect 2320 2540 2420 2560
rect 2460 2540 2560 2560
rect 2600 2540 2700 2560
rect 2740 2540 2840 2560
rect 2880 2540 2980 2560
rect 3020 2540 3120 2560
rect 3160 2540 3260 2560
rect 3300 2540 3400 2560
rect 3440 2540 3540 2560
rect 2180 2460 2280 2480
rect 2320 2460 2420 2480
rect 2460 2460 2560 2480
rect 2600 2460 2700 2480
rect 2740 2460 2840 2480
rect 2880 2460 2980 2480
rect 3020 2460 3120 2480
rect 3160 2460 3260 2480
rect 3300 2460 3400 2480
rect 3440 2460 3540 2480
rect -160 2350 -60 2360
rect -200 2340 -60 2350
rect -20 2350 80 2360
rect 120 2350 220 2360
rect -20 2340 220 2350
rect 260 2350 360 2360
rect 400 2350 500 2360
rect 260 2340 500 2350
rect 540 2350 640 2360
rect 680 2350 780 2360
rect 540 2340 780 2350
rect 820 2350 920 2360
rect 960 2350 1060 2360
rect 820 2340 1060 2350
rect 1100 2350 1200 2360
rect 1240 2350 1340 2360
rect 2040 2350 2140 2360
rect 2180 2350 2280 2360
rect 1100 2340 1340 2350
rect 1610 2340 1660 2350
rect -200 2320 -190 2340
rect -170 2330 -140 2340
rect 60 2330 90 2340
rect -170 2320 -160 2330
rect -200 2310 -160 2320
rect 80 2320 90 2330
rect 110 2330 140 2340
rect 340 2330 370 2340
rect 110 2320 120 2330
rect 80 2310 120 2320
rect 360 2320 370 2330
rect 390 2330 420 2340
rect 620 2330 650 2340
rect 390 2320 400 2330
rect 360 2310 400 2320
rect 640 2320 650 2330
rect 670 2330 700 2340
rect 900 2330 930 2340
rect 670 2320 680 2330
rect 640 2310 680 2320
rect 920 2320 930 2330
rect 950 2330 980 2340
rect 1180 2330 1210 2340
rect 950 2320 960 2330
rect 920 2310 960 2320
rect 1200 2320 1210 2330
rect 1230 2330 1260 2340
rect 1230 2320 1240 2330
rect 1200 2310 1240 2320
rect 1610 2320 1620 2340
rect 1640 2320 1660 2340
rect 1610 2310 1660 2320
rect 1640 2250 1660 2310
rect -90 2170 -50 2180
rect -90 2150 -80 2170
rect -60 2150 -50 2170
rect -20 2150 0 2250
rect 100 2210 120 2250
rect 150 2210 170 2250
rect 100 2190 170 2210
rect 100 2150 120 2190
rect 150 2150 170 2190
rect 270 2210 290 2250
rect 320 2210 340 2250
rect 270 2190 340 2210
rect 270 2150 290 2190
rect 320 2150 340 2190
rect 440 2210 460 2250
rect 490 2210 510 2250
rect 440 2190 510 2210
rect 440 2150 460 2190
rect 490 2150 510 2190
rect 610 2210 630 2250
rect 660 2210 680 2250
rect 610 2190 680 2210
rect 610 2150 630 2190
rect 660 2150 680 2190
rect 780 2210 800 2250
rect 830 2210 850 2250
rect 780 2190 850 2210
rect 780 2150 800 2190
rect 830 2150 850 2190
rect 950 2210 970 2250
rect 1000 2210 1020 2250
rect 950 2190 1020 2210
rect 950 2150 970 2190
rect 1000 2150 1020 2190
rect 1120 2210 1140 2250
rect 1170 2210 1190 2250
rect 1120 2190 1190 2210
rect 1120 2150 1140 2190
rect 1170 2150 1190 2190
rect 1290 2210 1310 2250
rect 1340 2210 1360 2250
rect 1290 2190 1360 2210
rect 1290 2150 1310 2190
rect 1340 2150 1360 2190
rect 1460 2210 1480 2250
rect 1510 2210 1530 2250
rect 1460 2190 1530 2210
rect 1460 2150 1480 2190
rect 1510 2150 1530 2190
rect 1630 2210 1660 2250
rect 1720 2340 1770 2350
rect 2040 2340 2280 2350
rect 2320 2350 2420 2360
rect 2460 2350 2560 2360
rect 2320 2340 2560 2350
rect 2600 2350 2700 2360
rect 2740 2350 2840 2360
rect 2600 2340 2840 2350
rect 2880 2350 2980 2360
rect 3020 2350 3120 2360
rect 2880 2340 3120 2350
rect 3160 2350 3260 2360
rect 3300 2350 3400 2360
rect 3160 2340 3400 2350
rect 3440 2350 3540 2360
rect 3440 2340 3580 2350
rect 1720 2320 1740 2340
rect 1760 2320 1770 2340
rect 2120 2330 2150 2340
rect 1720 2310 1770 2320
rect 2140 2320 2150 2330
rect 2170 2330 2200 2340
rect 2400 2330 2430 2340
rect 2170 2320 2180 2330
rect 2140 2310 2180 2320
rect 2420 2320 2430 2330
rect 2450 2330 2480 2340
rect 2680 2330 2710 2340
rect 2450 2320 2460 2330
rect 2420 2310 2460 2320
rect 2700 2320 2710 2330
rect 2730 2330 2760 2340
rect 2960 2330 2990 2340
rect 2730 2320 2740 2330
rect 2700 2310 2740 2320
rect 2980 2320 2990 2330
rect 3010 2330 3040 2340
rect 3240 2330 3270 2340
rect 3010 2320 3020 2330
rect 2980 2310 3020 2320
rect 3260 2320 3270 2330
rect 3290 2330 3320 2340
rect 3520 2330 3550 2340
rect 3290 2320 3300 2330
rect 3260 2310 3300 2320
rect 3540 2320 3550 2330
rect 3570 2320 3580 2340
rect 3540 2310 3580 2320
rect 1720 2250 1740 2310
rect 1720 2210 1750 2250
rect 1630 2190 1750 2210
rect 1630 2150 1650 2190
rect -90 2140 -50 2150
rect -70 2080 -50 2140
rect -300 1580 -280 2080
rect -80 2060 -50 2080
rect -80 1580 -60 2060
rect -300 1060 -280 1540
rect -310 1040 -280 1060
rect -80 1040 -60 1540
rect -20 1040 0 2040
rect 100 1550 120 2040
rect 150 1550 170 2040
rect 100 1530 170 1550
rect 100 1040 120 1530
rect 150 1040 170 1530
rect 270 1550 290 2040
rect 320 1550 340 2040
rect 270 1530 340 1550
rect 270 1040 290 1530
rect 320 1040 340 1530
rect 440 1550 460 2040
rect 490 1550 510 2040
rect 440 1530 510 1550
rect 440 1040 460 1530
rect 490 1040 510 1530
rect 610 1550 630 2040
rect 660 1550 680 2040
rect 610 1530 680 1550
rect 610 1040 630 1530
rect 660 1040 680 1530
rect 780 1550 800 2040
rect 830 1550 850 2040
rect 780 1530 850 1550
rect 780 1040 800 1530
rect 830 1040 850 1530
rect 950 1550 970 2040
rect 1000 1550 1020 2040
rect 950 1530 1020 1550
rect 950 1040 970 1530
rect 1000 1040 1020 1530
rect 1120 1550 1140 2040
rect 1170 1550 1190 2040
rect 1120 1530 1190 1550
rect 1120 1040 1140 1530
rect 1170 1040 1190 1530
rect 1290 1550 1310 2040
rect 1340 1550 1360 2040
rect 1290 1530 1360 1550
rect 1290 1040 1310 1530
rect 1340 1040 1360 1530
rect 1460 1550 1480 2040
rect 1510 1550 1530 2040
rect 1460 1530 1530 1550
rect 1460 1040 1480 1530
rect 1510 1040 1530 1530
rect 1630 1550 1650 2040
rect 1680 1550 1700 2190
rect 1730 2150 1750 2190
rect 1850 2210 1870 2250
rect 1900 2210 1920 2250
rect 1850 2190 1920 2210
rect 1850 2150 1870 2190
rect 1900 2150 1920 2190
rect 2020 2210 2040 2250
rect 2070 2210 2090 2250
rect 2020 2190 2090 2210
rect 2020 2150 2040 2190
rect 2070 2150 2090 2190
rect 2190 2210 2210 2250
rect 2240 2210 2260 2250
rect 2190 2190 2260 2210
rect 2190 2150 2210 2190
rect 2240 2150 2260 2190
rect 2360 2210 2380 2250
rect 2410 2210 2430 2250
rect 2360 2190 2430 2210
rect 2360 2150 2380 2190
rect 2410 2150 2430 2190
rect 2530 2210 2550 2250
rect 2580 2210 2600 2250
rect 2530 2190 2600 2210
rect 2530 2150 2550 2190
rect 2580 2150 2600 2190
rect 2700 2210 2720 2250
rect 2750 2210 2770 2250
rect 2700 2190 2770 2210
rect 2700 2150 2720 2190
rect 2750 2150 2770 2190
rect 2870 2210 2890 2250
rect 2920 2210 2940 2250
rect 2870 2190 2940 2210
rect 2870 2150 2890 2190
rect 2920 2150 2940 2190
rect 3040 2210 3060 2250
rect 3090 2210 3110 2250
rect 3040 2190 3110 2210
rect 3040 2150 3060 2190
rect 3090 2150 3110 2190
rect 3210 2210 3230 2250
rect 3260 2210 3280 2250
rect 3210 2190 3280 2210
rect 3210 2150 3230 2190
rect 3260 2150 3280 2190
rect 3380 2150 3400 2250
rect 3430 2170 3470 2180
rect 3430 2150 3440 2170
rect 3460 2150 3470 2170
rect 3430 2140 3470 2150
rect 3430 2080 3450 2140
rect 3430 2060 3460 2080
rect 1730 1550 1750 2040
rect 1630 1530 1750 1550
rect 1630 1040 1650 1530
rect 1730 1040 1750 1530
rect 1850 1550 1870 2040
rect 1900 1550 1920 2040
rect 1850 1530 1920 1550
rect 1850 1040 1870 1530
rect 1900 1040 1920 1530
rect 2020 1550 2040 2040
rect 2070 1550 2090 2040
rect 2020 1530 2090 1550
rect 2020 1040 2040 1530
rect 2070 1040 2090 1530
rect 2190 1550 2210 2040
rect 2240 1550 2260 2040
rect 2190 1530 2260 1550
rect 2190 1040 2210 1530
rect 2240 1040 2260 1530
rect 2360 1550 2380 2040
rect 2410 1550 2430 2040
rect 2360 1530 2430 1550
rect 2360 1040 2380 1530
rect 2410 1040 2430 1530
rect 2530 1550 2550 2040
rect 2580 1550 2600 2040
rect 2530 1530 2600 1550
rect 2530 1040 2550 1530
rect 2580 1040 2600 1530
rect 2700 1550 2720 2040
rect 2750 1550 2770 2040
rect 2700 1530 2770 1550
rect 2700 1040 2720 1530
rect 2750 1040 2770 1530
rect 2870 1550 2890 2040
rect 2920 1550 2940 2040
rect 2870 1530 2940 1550
rect 2870 1040 2890 1530
rect 2920 1040 2940 1530
rect 3040 1550 3060 2040
rect 3090 1550 3110 2040
rect 3040 1530 3110 1550
rect 3040 1040 3060 1530
rect 3090 1040 3110 1530
rect 3210 1550 3230 2040
rect 3260 1550 3280 2040
rect 3210 1530 3280 1550
rect 3210 1040 3230 1530
rect 3260 1040 3280 1530
rect 3380 1040 3400 2040
rect 3440 1580 3460 2060
rect 3660 1580 3680 2080
rect 3440 1040 3460 1540
rect 3660 1060 3680 1540
rect 3660 1040 3690 1060
rect -310 980 -290 1040
rect -310 970 -270 980
rect -310 950 -300 970
rect -280 950 -270 970
rect -310 940 -270 950
rect -20 20 0 1000
rect -40 0 0 20
rect 100 510 120 1000
rect 150 510 170 1000
rect 100 490 170 510
rect 100 0 120 490
rect 150 0 170 490
rect 270 510 290 1000
rect 320 510 340 1000
rect 270 490 340 510
rect 270 0 290 490
rect 320 0 340 490
rect 440 510 460 1000
rect 490 510 510 1000
rect 440 490 510 510
rect 440 0 460 490
rect 490 0 510 490
rect 610 510 630 1000
rect 660 510 680 1000
rect 610 490 680 510
rect 610 0 630 490
rect 660 0 680 490
rect 780 510 800 1000
rect 830 510 850 1000
rect 780 490 850 510
rect 780 0 800 490
rect 830 0 850 490
rect 950 510 970 1000
rect 1000 510 1020 1000
rect 950 490 1020 510
rect 950 0 970 490
rect 1000 0 1020 490
rect 1120 510 1140 1000
rect 1170 510 1190 1000
rect 1120 490 1190 510
rect 1120 0 1140 490
rect 1170 0 1190 490
rect 1290 510 1310 1000
rect 1340 510 1360 1000
rect 1290 490 1360 510
rect 1290 0 1310 490
rect 1340 0 1360 490
rect 1460 510 1480 1000
rect 1510 510 1530 1000
rect 1460 490 1530 510
rect 1460 0 1480 490
rect 1510 0 1530 490
rect 1630 510 1650 1000
rect 1730 510 1750 1000
rect 1630 490 1750 510
rect 1630 0 1650 490
rect 1730 0 1750 490
rect 1850 510 1870 1000
rect 1900 510 1920 1000
rect 1850 490 1920 510
rect 1850 0 1870 490
rect 1900 0 1920 490
rect 2020 510 2040 1000
rect 2070 510 2090 1000
rect 2020 490 2090 510
rect 2020 0 2040 490
rect 2070 0 2090 490
rect 2190 510 2210 1000
rect 2240 510 2260 1000
rect 2190 490 2260 510
rect 2190 0 2210 490
rect 2240 0 2260 490
rect 2360 510 2380 1000
rect 2410 510 2430 1000
rect 2360 490 2430 510
rect 2360 0 2380 490
rect 2410 0 2430 490
rect 2530 510 2550 1000
rect 2580 510 2600 1000
rect 2530 490 2600 510
rect 2530 0 2550 490
rect 2580 0 2600 490
rect 2700 510 2720 1000
rect 2750 510 2770 1000
rect 2700 490 2770 510
rect 2700 0 2720 490
rect 2750 0 2770 490
rect 2870 510 2890 1000
rect 2920 510 2940 1000
rect 2870 490 2940 510
rect 2870 0 2890 490
rect 2920 0 2940 490
rect 3040 510 3060 1000
rect 3090 510 3110 1000
rect 3040 490 3110 510
rect 3040 0 3060 490
rect 3090 0 3110 490
rect 3210 510 3230 1000
rect 3260 510 3280 1000
rect 3210 490 3280 510
rect 3210 0 3230 490
rect 3260 0 3280 490
rect 3380 20 3400 1000
rect 3670 980 3690 1040
rect 3650 970 3690 980
rect 3650 950 3660 970
rect 3680 950 3690 970
rect 3650 940 3690 950
rect 3380 0 3420 20
rect -40 -20 -20 0
rect -60 -30 -20 -20
rect -60 -50 -50 -30
rect -30 -50 -20 -30
rect -60 -60 -20 -50
rect 3400 -20 3420 0
rect 3400 -30 3440 -20
rect 3400 -50 3410 -30
rect 3430 -50 3440 -30
rect 3400 -60 3440 -50
<< polycont >>
rect -50 5050 -30 5070
rect 3410 5050 3430 5070
rect -300 4050 -280 4070
rect 3660 4050 3680 4070
rect -80 2850 -60 2870
rect -190 2680 -170 2700
rect 90 2680 110 2700
rect 370 2680 390 2700
rect 650 2680 670 2700
rect 930 2680 950 2700
rect 1210 2680 1230 2700
rect 1620 2680 1640 2700
rect 3440 2850 3460 2870
rect 1740 2680 1760 2700
rect 2150 2680 2170 2700
rect 2430 2680 2450 2700
rect 2710 2680 2730 2700
rect 2990 2680 3010 2700
rect 3270 2680 3290 2700
rect 3550 2680 3570 2700
rect -190 2320 -170 2340
rect 90 2320 110 2340
rect 370 2320 390 2340
rect 650 2320 670 2340
rect 930 2320 950 2340
rect 1210 2320 1230 2340
rect 1620 2320 1640 2340
rect -80 2150 -60 2170
rect 1740 2320 1760 2340
rect 2150 2320 2170 2340
rect 2430 2320 2450 2340
rect 2710 2320 2730 2340
rect 2990 2320 3010 2340
rect 3270 2320 3290 2340
rect 3550 2320 3570 2340
rect 3440 2150 3460 2170
rect -300 950 -280 970
rect 3660 950 3680 970
rect -50 -50 -30 -30
rect 3410 -50 3430 -30
<< locali >>
rect -60 5070 -20 5080
rect 20 5070 30 5090
rect 70 5070 80 5090
rect 190 5070 200 5090
rect 240 5070 250 5090
rect 360 5070 370 5090
rect 410 5070 420 5090
rect 530 5070 540 5090
rect 580 5070 590 5090
rect 700 5070 710 5090
rect 750 5070 760 5090
rect 870 5070 880 5090
rect 920 5070 930 5090
rect 1040 5070 1050 5090
rect 1090 5070 1100 5090
rect 1210 5070 1220 5090
rect 1260 5070 1270 5090
rect 1380 5070 1390 5090
rect 1430 5070 1440 5090
rect 1550 5070 1560 5090
rect 1600 5070 1610 5090
rect 1770 5070 1780 5090
rect 1820 5070 1830 5090
rect 1940 5070 1950 5090
rect 1990 5070 2000 5090
rect 2110 5070 2120 5090
rect 2160 5070 2170 5090
rect 2280 5070 2290 5090
rect 2330 5070 2340 5090
rect 2450 5070 2460 5090
rect 2500 5070 2510 5090
rect 2620 5070 2630 5090
rect 2670 5070 2680 5090
rect 2790 5070 2800 5090
rect 2840 5070 2850 5090
rect 2960 5070 2970 5090
rect 3010 5070 3020 5090
rect 3130 5070 3140 5090
rect 3180 5070 3190 5090
rect 3300 5070 3310 5090
rect 3350 5070 3360 5090
rect 3400 5070 3440 5080
rect -60 5050 -50 5070
rect -30 5050 3410 5070
rect 3430 5050 3440 5070
rect -60 5040 -20 5050
rect 20 5030 30 5050
rect 70 5030 80 5050
rect 20 5020 80 5030
rect 190 5030 200 5050
rect 240 5030 250 5050
rect 190 5020 250 5030
rect 360 5030 370 5050
rect 410 5030 420 5050
rect 360 5020 420 5030
rect 530 5030 540 5050
rect 580 5030 590 5050
rect 530 5020 590 5030
rect 700 5030 710 5050
rect 750 5030 760 5050
rect 700 5020 760 5030
rect 870 5030 880 5050
rect 920 5030 930 5050
rect 870 5020 930 5030
rect 1040 5030 1050 5050
rect 1090 5030 1100 5050
rect 1040 5020 1100 5030
rect 1210 5030 1220 5050
rect 1260 5030 1270 5050
rect 1210 5020 1270 5030
rect 1380 5030 1390 5050
rect 1430 5030 1440 5050
rect 1380 5020 1440 5030
rect 1550 5030 1560 5050
rect 1600 5030 1610 5050
rect 1550 5020 1610 5030
rect -310 4070 -270 4080
rect -310 4050 -300 4070
rect -280 4050 -170 4070
rect -310 4040 -270 4050
rect -190 4020 -170 4050
rect -210 4010 -150 4020
rect -210 3990 -200 4010
rect -160 3990 -150 4010
rect -210 3980 -150 3990
rect 20 4010 80 4020
rect 20 3990 30 4010
rect 70 3990 80 4010
rect 20 3980 80 3990
rect 190 4010 250 4020
rect 190 3990 200 4010
rect 240 3990 250 4010
rect 190 3980 250 3990
rect 360 4010 420 4020
rect 360 3990 370 4010
rect 410 3990 420 4010
rect 360 3980 420 3990
rect 530 4010 590 4020
rect 530 3990 540 4010
rect 580 3990 590 4010
rect 530 3980 590 3990
rect 700 4010 760 4020
rect 700 3990 710 4010
rect 750 3990 760 4010
rect 700 3980 760 3990
rect 870 4010 930 4020
rect 870 3990 880 4010
rect 920 3990 930 4010
rect 870 3980 930 3990
rect 1040 4010 1100 4020
rect 1040 3990 1050 4010
rect 1090 3990 1100 4010
rect 1040 3980 1100 3990
rect 1210 4010 1270 4020
rect 1210 3990 1220 4010
rect 1260 3990 1270 4010
rect 1210 3980 1270 3990
rect 1380 4010 1440 4020
rect 1380 3990 1390 4010
rect 1430 3990 1440 4010
rect 1380 3980 1440 3990
rect 1550 4010 1610 4020
rect 1550 3990 1560 4010
rect 1600 3990 1610 4010
rect 1550 3980 1610 3990
rect -210 3470 -150 3480
rect -210 3450 -200 3470
rect -160 3450 -110 3470
rect -210 3440 -150 3450
rect -210 2930 -150 2940
rect -210 2910 -200 2930
rect -160 2910 -150 2930
rect -210 2900 -150 2910
rect -190 2710 -170 2900
rect -130 2720 -110 3450
rect 20 2970 80 2980
rect 20 2950 30 2970
rect 70 2950 80 2970
rect 190 2970 250 2980
rect 190 2950 200 2970
rect 240 2950 250 2970
rect 360 2970 420 2980
rect 360 2950 370 2970
rect 410 2950 420 2970
rect 530 2970 590 2980
rect 530 2950 540 2970
rect 580 2950 590 2970
rect 700 2970 760 2980
rect 700 2950 710 2970
rect 750 2950 760 2970
rect 870 2970 930 2980
rect 870 2950 880 2970
rect 920 2950 930 2970
rect 1040 2970 1100 2980
rect 1040 2950 1050 2970
rect 1090 2950 1100 2970
rect 1210 2970 1270 2980
rect 1210 2950 1220 2970
rect 1260 2950 1270 2970
rect 1380 2970 1440 2980
rect 1380 2950 1390 2970
rect 1430 2950 1440 2970
rect 1550 2970 1610 2980
rect 1550 2950 1560 2970
rect 1600 2950 1610 2970
rect 1680 2950 1700 5050
rect 1770 5030 1780 5050
rect 1820 5030 1830 5050
rect 1770 5020 1830 5030
rect 1940 5030 1950 5050
rect 1990 5030 2000 5050
rect 1940 5020 2000 5030
rect 2110 5030 2120 5050
rect 2160 5030 2170 5050
rect 2110 5020 2170 5030
rect 2280 5030 2290 5050
rect 2330 5030 2340 5050
rect 2280 5020 2340 5030
rect 2450 5030 2460 5050
rect 2500 5030 2510 5050
rect 2450 5020 2510 5030
rect 2620 5030 2630 5050
rect 2670 5030 2680 5050
rect 2620 5020 2680 5030
rect 2790 5030 2800 5050
rect 2840 5030 2850 5050
rect 2790 5020 2850 5030
rect 2960 5030 2970 5050
rect 3010 5030 3020 5050
rect 2960 5020 3020 5030
rect 3130 5030 3140 5050
rect 3180 5030 3190 5050
rect 3130 5020 3190 5030
rect 3300 5030 3310 5050
rect 3350 5030 3360 5050
rect 3400 5040 3440 5050
rect 3300 5020 3360 5030
rect 3650 4070 3690 4080
rect 3550 4050 3660 4070
rect 3680 4050 3690 4070
rect 3550 4020 3570 4050
rect 3650 4040 3690 4050
rect 1770 4010 1830 4020
rect 1770 3990 1780 4010
rect 1820 3990 1830 4010
rect 1770 3980 1830 3990
rect 1940 4010 2000 4020
rect 1940 3990 1950 4010
rect 1990 3990 2000 4010
rect 1940 3980 2000 3990
rect 2110 4010 2170 4020
rect 2110 3990 2120 4010
rect 2160 3990 2170 4010
rect 2110 3980 2170 3990
rect 2280 4010 2340 4020
rect 2280 3990 2290 4010
rect 2330 3990 2340 4010
rect 2280 3980 2340 3990
rect 2450 4010 2510 4020
rect 2450 3990 2460 4010
rect 2500 3990 2510 4010
rect 2450 3980 2510 3990
rect 2620 4010 2680 4020
rect 2620 3990 2630 4010
rect 2670 3990 2680 4010
rect 2620 3980 2680 3990
rect 2790 4010 2850 4020
rect 2790 3990 2800 4010
rect 2840 3990 2850 4010
rect 2790 3980 2850 3990
rect 2960 4010 3020 4020
rect 2960 3990 2970 4010
rect 3010 3990 3020 4010
rect 2960 3980 3020 3990
rect 3130 4010 3190 4020
rect 3130 3990 3140 4010
rect 3180 3990 3190 4010
rect 3130 3980 3190 3990
rect 3300 4010 3360 4020
rect 3300 3990 3310 4010
rect 3350 3990 3360 4010
rect 3300 3980 3360 3990
rect 3530 4010 3590 4020
rect 3530 3990 3540 4010
rect 3580 3990 3590 4010
rect 3530 3980 3590 3990
rect 3530 3470 3590 3480
rect 3490 3450 3540 3470
rect 3580 3450 3590 3470
rect 1770 2970 1830 2980
rect 1770 2950 1780 2970
rect 1820 2950 1830 2970
rect 1940 2970 2000 2980
rect 1940 2950 1950 2970
rect 1990 2950 2000 2970
rect 2110 2970 2170 2980
rect 2110 2950 2120 2970
rect 2160 2950 2170 2970
rect 2280 2970 2340 2980
rect 2280 2950 2290 2970
rect 2330 2950 2340 2970
rect 2450 2970 2510 2980
rect 2450 2950 2460 2970
rect 2500 2950 2510 2970
rect 2620 2970 2680 2980
rect 2620 2950 2630 2970
rect 2670 2950 2680 2970
rect 2790 2970 2850 2980
rect 2790 2950 2800 2970
rect 2840 2950 2850 2970
rect 2960 2970 3020 2980
rect 2960 2950 2970 2970
rect 3010 2950 3020 2970
rect 3130 2970 3190 2980
rect 3130 2950 3140 2970
rect 3180 2950 3190 2970
rect 3300 2970 3360 2980
rect 3300 2950 3310 2970
rect 3350 2950 3360 2970
rect 20 2930 3360 2950
rect 20 2910 30 2930
rect 70 2910 80 2930
rect 20 2900 80 2910
rect 190 2910 200 2930
rect 240 2910 250 2930
rect 190 2900 250 2910
rect 360 2910 370 2930
rect 410 2910 420 2930
rect 360 2900 420 2910
rect 530 2910 540 2930
rect 580 2910 590 2930
rect 530 2900 590 2910
rect 700 2910 710 2930
rect 750 2910 760 2930
rect 700 2900 760 2910
rect 870 2910 880 2930
rect 920 2910 930 2930
rect 870 2900 930 2910
rect 1040 2910 1050 2930
rect 1090 2910 1100 2930
rect 1040 2900 1100 2910
rect 1210 2910 1220 2930
rect 1260 2910 1270 2930
rect 1210 2900 1270 2910
rect 1380 2910 1390 2930
rect 1430 2910 1440 2930
rect 1380 2900 1440 2910
rect 1550 2910 1560 2930
rect 1600 2910 1610 2930
rect 1550 2900 1610 2910
rect -90 2870 -50 2880
rect -90 2850 -80 2870
rect -60 2850 -50 2870
rect -90 2840 -50 2850
rect -80 2760 -60 2840
rect 20 2760 80 2770
rect 190 2760 250 2770
rect 360 2760 420 2770
rect 530 2760 590 2770
rect 700 2760 760 2770
rect 870 2760 930 2770
rect 1040 2760 1100 2770
rect 1210 2760 1270 2770
rect 1380 2760 1440 2770
rect 1550 2760 1610 2770
rect -80 2740 30 2760
rect 70 2740 200 2760
rect 240 2740 370 2760
rect 410 2740 540 2760
rect 580 2740 710 2760
rect 750 2740 880 2760
rect 920 2740 1050 2760
rect 1090 2740 1220 2760
rect 1260 2740 1390 2760
rect 1430 2740 1560 2760
rect 1600 2740 1610 2760
rect 20 2730 80 2740
rect 190 2730 250 2740
rect 360 2730 420 2740
rect 530 2730 590 2740
rect 700 2730 760 2740
rect 870 2730 930 2740
rect 1040 2730 1100 2740
rect 1210 2730 1270 2740
rect 1380 2730 1440 2740
rect 1550 2730 1610 2740
rect -200 2700 -160 2710
rect -130 2700 -30 2720
rect -200 2680 -190 2700
rect -170 2680 -160 2700
rect -200 2670 -160 2680
rect -190 2640 -170 2670
rect -50 2640 -30 2700
rect 80 2700 120 2710
rect 360 2700 400 2710
rect 640 2700 680 2710
rect 920 2700 960 2710
rect 1200 2700 1240 2710
rect 1550 2700 1570 2730
rect 80 2680 90 2700
rect 110 2680 370 2700
rect 390 2680 650 2700
rect 670 2680 930 2700
rect 950 2680 1210 2700
rect 1230 2680 1570 2700
rect 80 2670 120 2680
rect 360 2670 400 2680
rect 640 2670 680 2680
rect 920 2670 960 2680
rect 1200 2670 1240 2680
rect 1550 2670 1570 2680
rect 1610 2700 1650 2710
rect 1610 2680 1620 2700
rect 1640 2680 1650 2700
rect 1610 2670 1650 2680
rect 90 2640 110 2670
rect 370 2640 390 2670
rect 650 2640 670 2670
rect 930 2640 950 2670
rect 1210 2640 1230 2670
rect 1550 2660 1590 2670
rect 1550 2640 1560 2660
rect 1580 2640 1590 2660
rect -240 2630 -160 2640
rect -240 2590 -230 2630
rect -210 2590 -190 2630
rect -170 2590 -160 2630
rect -240 2580 -160 2590
rect -60 2630 -20 2640
rect -60 2590 -50 2630
rect -30 2590 -20 2630
rect -60 2580 -20 2590
rect 80 2630 120 2640
rect 80 2590 90 2630
rect 110 2590 120 2630
rect 80 2580 120 2590
rect 220 2630 260 2640
rect 220 2590 230 2630
rect 250 2590 260 2630
rect 220 2580 260 2590
rect 360 2630 400 2640
rect 360 2590 370 2630
rect 390 2590 400 2630
rect 360 2580 400 2590
rect 500 2630 540 2640
rect 500 2590 510 2630
rect 530 2590 540 2630
rect 500 2580 540 2590
rect 640 2630 680 2640
rect 640 2590 650 2630
rect 670 2590 680 2630
rect 640 2580 680 2590
rect 780 2630 820 2640
rect 780 2590 790 2630
rect 810 2590 820 2630
rect 780 2580 820 2590
rect 920 2630 960 2640
rect 920 2590 930 2630
rect 950 2590 960 2630
rect 920 2580 960 2590
rect 1060 2630 1100 2640
rect 1060 2590 1070 2630
rect 1090 2590 1100 2630
rect 1060 2580 1100 2590
rect 1200 2630 1240 2640
rect 1200 2590 1210 2630
rect 1230 2590 1240 2630
rect 1200 2580 1240 2590
rect 1340 2630 1380 2640
rect 1550 2630 1590 2640
rect 1340 2590 1350 2630
rect 1370 2600 1380 2630
rect 1370 2590 1590 2600
rect 1340 2580 1560 2590
rect -190 2520 -170 2580
rect -50 2560 -30 2580
rect 230 2560 250 2580
rect 510 2560 530 2580
rect 790 2560 810 2580
rect 1070 2560 1090 2580
rect 1350 2560 1370 2580
rect 1550 2570 1560 2580
rect 1580 2570 1590 2590
rect 1550 2560 1590 2570
rect -50 2540 1370 2560
rect 1410 2520 1450 2530
rect 1550 2520 1590 2530
rect -190 2500 1420 2520
rect 1440 2500 1560 2520
rect 1580 2500 1590 2520
rect -190 2440 -170 2500
rect 1410 2490 1450 2500
rect 1550 2490 1590 2500
rect -50 2460 1370 2480
rect -50 2440 -30 2460
rect 230 2440 250 2460
rect 510 2440 530 2460
rect 790 2440 810 2460
rect 1070 2440 1090 2460
rect 1350 2440 1370 2460
rect 1550 2450 1590 2460
rect 1550 2440 1560 2450
rect -240 2430 -160 2440
rect -240 2390 -230 2430
rect -210 2390 -190 2430
rect -170 2390 -160 2430
rect -240 2380 -160 2390
rect -60 2430 -20 2440
rect -60 2390 -50 2430
rect -30 2390 -20 2430
rect -60 2380 -20 2390
rect 80 2430 120 2440
rect 80 2390 90 2430
rect 110 2390 120 2430
rect 80 2380 120 2390
rect 220 2430 260 2440
rect 220 2390 230 2430
rect 250 2390 260 2430
rect 220 2380 260 2390
rect 360 2430 400 2440
rect 360 2390 370 2430
rect 390 2390 400 2430
rect 360 2380 400 2390
rect 500 2430 540 2440
rect 500 2390 510 2430
rect 530 2390 540 2430
rect 500 2380 540 2390
rect 640 2430 680 2440
rect 640 2390 650 2430
rect 670 2390 680 2430
rect 640 2380 680 2390
rect 780 2430 820 2440
rect 780 2390 790 2430
rect 810 2390 820 2430
rect 780 2380 820 2390
rect 920 2430 960 2440
rect 920 2390 930 2430
rect 950 2390 960 2430
rect 920 2380 960 2390
rect 1060 2430 1100 2440
rect 1060 2390 1070 2430
rect 1090 2390 1100 2430
rect 1060 2380 1100 2390
rect 1200 2430 1240 2440
rect 1200 2390 1210 2430
rect 1230 2390 1240 2430
rect 1200 2380 1240 2390
rect 1340 2430 1560 2440
rect 1580 2430 1590 2450
rect 1340 2390 1350 2430
rect 1370 2420 1590 2430
rect 1370 2390 1380 2420
rect 1340 2380 1380 2390
rect 1550 2380 1590 2390
rect -190 2350 -170 2380
rect -200 2340 -160 2350
rect -200 2320 -190 2340
rect -170 2320 -160 2340
rect -50 2320 -30 2380
rect 90 2350 110 2380
rect 370 2350 390 2380
rect 650 2350 670 2380
rect 930 2350 950 2380
rect 1210 2350 1230 2380
rect 1550 2360 1560 2380
rect 1580 2360 1590 2380
rect 1550 2350 1590 2360
rect 1620 2350 1640 2670
rect -200 2310 -160 2320
rect -190 2120 -170 2310
rect -130 2300 -30 2320
rect 80 2340 120 2350
rect 360 2340 400 2350
rect 640 2340 680 2350
rect 920 2340 960 2350
rect 1200 2340 1240 2350
rect 1550 2340 1570 2350
rect 80 2320 90 2340
rect 110 2320 370 2340
rect 390 2320 650 2340
rect 670 2320 930 2340
rect 950 2320 1210 2340
rect 1230 2320 1570 2340
rect 80 2310 120 2320
rect 360 2310 400 2320
rect 640 2310 680 2320
rect 920 2310 960 2320
rect 1200 2310 1240 2320
rect -210 2110 -150 2120
rect -210 2090 -200 2110
rect -160 2090 -150 2110
rect -210 2080 -150 2090
rect -210 1570 -150 1580
rect -130 1570 -110 2300
rect 1550 2290 1570 2320
rect 1610 2340 1650 2350
rect 1610 2320 1620 2340
rect 1640 2320 1650 2340
rect 1610 2310 1650 2320
rect 20 2280 80 2290
rect 190 2280 250 2290
rect 360 2280 420 2290
rect 530 2280 590 2290
rect 700 2280 760 2290
rect 870 2280 930 2290
rect 1040 2280 1100 2290
rect 1210 2280 1270 2290
rect 1380 2280 1440 2290
rect 1550 2280 1610 2290
rect -80 2260 30 2280
rect 70 2260 200 2280
rect 240 2260 370 2280
rect 410 2260 540 2280
rect 580 2260 710 2280
rect 750 2260 880 2280
rect 920 2260 1050 2280
rect 1090 2260 1220 2280
rect 1260 2260 1390 2280
rect 1430 2260 1560 2280
rect 1600 2260 1610 2280
rect -80 2180 -60 2260
rect 20 2250 80 2260
rect 190 2250 250 2260
rect 360 2250 420 2260
rect 530 2250 590 2260
rect 700 2250 760 2260
rect 870 2250 930 2260
rect 1040 2250 1100 2260
rect 1210 2250 1270 2260
rect 1380 2250 1440 2260
rect 1550 2250 1610 2260
rect -90 2170 -50 2180
rect -90 2150 -80 2170
rect -60 2150 -50 2170
rect -90 2140 -50 2150
rect 20 2110 80 2120
rect 20 2090 30 2110
rect 70 2090 80 2110
rect 190 2110 250 2120
rect 190 2090 200 2110
rect 240 2090 250 2110
rect 360 2110 420 2120
rect 360 2090 370 2110
rect 410 2090 420 2110
rect 530 2110 590 2120
rect 530 2090 540 2110
rect 580 2090 590 2110
rect 700 2110 760 2120
rect 700 2090 710 2110
rect 750 2090 760 2110
rect 870 2110 930 2120
rect 870 2090 880 2110
rect 920 2090 930 2110
rect 1040 2110 1100 2120
rect 1040 2090 1050 2110
rect 1090 2090 1100 2110
rect 1210 2110 1270 2120
rect 1210 2090 1220 2110
rect 1260 2090 1270 2110
rect 1380 2110 1440 2120
rect 1380 2090 1390 2110
rect 1430 2090 1440 2110
rect 1550 2110 1610 2120
rect 1550 2090 1560 2110
rect 1600 2090 1610 2110
rect 1680 2090 1700 2930
rect 1770 2910 1780 2930
rect 1820 2910 1830 2930
rect 1770 2900 1830 2910
rect 1940 2910 1950 2930
rect 1990 2910 2000 2930
rect 1940 2900 2000 2910
rect 2110 2910 2120 2930
rect 2160 2910 2170 2930
rect 2110 2900 2170 2910
rect 2280 2910 2290 2930
rect 2330 2910 2340 2930
rect 2280 2900 2340 2910
rect 2450 2910 2460 2930
rect 2500 2910 2510 2930
rect 2450 2900 2510 2910
rect 2620 2910 2630 2930
rect 2670 2910 2680 2930
rect 2620 2900 2680 2910
rect 2790 2910 2800 2930
rect 2840 2910 2850 2930
rect 2790 2900 2850 2910
rect 2960 2910 2970 2930
rect 3010 2910 3020 2930
rect 2960 2900 3020 2910
rect 3130 2910 3140 2930
rect 3180 2910 3190 2930
rect 3130 2900 3190 2910
rect 3300 2910 3310 2930
rect 3350 2910 3360 2930
rect 3300 2900 3360 2910
rect 3430 2870 3470 2880
rect 3430 2850 3440 2870
rect 3460 2850 3470 2870
rect 3430 2840 3470 2850
rect 1770 2760 1830 2770
rect 1940 2760 2000 2770
rect 2110 2760 2170 2770
rect 2280 2760 2340 2770
rect 2450 2760 2510 2770
rect 2620 2760 2680 2770
rect 2790 2760 2850 2770
rect 2960 2760 3020 2770
rect 3130 2760 3190 2770
rect 3300 2760 3360 2770
rect 3440 2760 3460 2840
rect 1770 2740 1780 2760
rect 1820 2740 1950 2760
rect 1990 2740 2120 2760
rect 2160 2740 2290 2760
rect 2330 2740 2460 2760
rect 2500 2740 2630 2760
rect 2670 2740 2800 2760
rect 2840 2740 2970 2760
rect 3010 2740 3140 2760
rect 3180 2740 3310 2760
rect 3350 2740 3460 2760
rect 1770 2730 1830 2740
rect 1940 2730 2000 2740
rect 2110 2730 2170 2740
rect 2280 2730 2340 2740
rect 2450 2730 2510 2740
rect 2620 2730 2680 2740
rect 2790 2730 2850 2740
rect 2960 2730 3020 2740
rect 3130 2730 3190 2740
rect 3300 2730 3360 2740
rect 1730 2700 1770 2710
rect 1730 2680 1740 2700
rect 1760 2680 1770 2700
rect 1730 2670 1770 2680
rect 1810 2700 1830 2730
rect 3490 2720 3510 3450
rect 3530 3440 3590 3450
rect 3530 2930 3590 2940
rect 3530 2910 3540 2930
rect 3580 2910 3590 2930
rect 3530 2900 3590 2910
rect 2140 2700 2180 2710
rect 2420 2700 2460 2710
rect 2700 2700 2740 2710
rect 2980 2700 3020 2710
rect 3260 2700 3300 2710
rect 1810 2680 2150 2700
rect 2170 2680 2430 2700
rect 2450 2680 2710 2700
rect 2730 2680 2990 2700
rect 3010 2680 3270 2700
rect 3290 2680 3300 2700
rect 1810 2670 1830 2680
rect 2140 2670 2180 2680
rect 2420 2670 2460 2680
rect 2700 2670 2740 2680
rect 2980 2670 3020 2680
rect 3260 2670 3300 2680
rect 3410 2700 3510 2720
rect 3550 2710 3570 2900
rect 3540 2700 3580 2710
rect 1740 2350 1760 2670
rect 1790 2660 1830 2670
rect 1790 2640 1800 2660
rect 1820 2640 1830 2660
rect 2150 2640 2170 2670
rect 2430 2640 2450 2670
rect 2710 2640 2730 2670
rect 2990 2640 3010 2670
rect 3270 2640 3290 2670
rect 3410 2640 3430 2700
rect 3540 2680 3550 2700
rect 3570 2680 3580 2700
rect 3540 2670 3580 2680
rect 3550 2640 3570 2670
rect 1790 2630 1830 2640
rect 2000 2630 2040 2640
rect 2000 2600 2010 2630
rect 1790 2590 2010 2600
rect 2030 2590 2040 2630
rect 1790 2570 1800 2590
rect 1820 2580 2040 2590
rect 2140 2630 2180 2640
rect 2140 2590 2150 2630
rect 2170 2590 2180 2630
rect 2140 2580 2180 2590
rect 2280 2630 2320 2640
rect 2280 2590 2290 2630
rect 2310 2590 2320 2630
rect 2280 2580 2320 2590
rect 2420 2630 2460 2640
rect 2420 2590 2430 2630
rect 2450 2590 2460 2630
rect 2420 2580 2460 2590
rect 2560 2630 2600 2640
rect 2560 2590 2570 2630
rect 2590 2590 2600 2630
rect 2560 2580 2600 2590
rect 2700 2630 2740 2640
rect 2700 2590 2710 2630
rect 2730 2590 2740 2630
rect 2700 2580 2740 2590
rect 2840 2630 2880 2640
rect 2840 2590 2850 2630
rect 2870 2590 2880 2630
rect 2840 2580 2880 2590
rect 2980 2630 3020 2640
rect 2980 2590 2990 2630
rect 3010 2590 3020 2630
rect 2980 2580 3020 2590
rect 3120 2630 3160 2640
rect 3120 2590 3130 2630
rect 3150 2590 3160 2630
rect 3120 2580 3160 2590
rect 3260 2630 3300 2640
rect 3260 2590 3270 2630
rect 3290 2590 3300 2630
rect 3260 2580 3300 2590
rect 3400 2630 3440 2640
rect 3400 2590 3410 2630
rect 3430 2590 3440 2630
rect 3400 2580 3440 2590
rect 3540 2630 3620 2640
rect 3540 2590 3550 2630
rect 3570 2590 3590 2630
rect 3610 2590 3620 2630
rect 3540 2580 3620 2590
rect 1820 2570 1830 2580
rect 1790 2560 1830 2570
rect 2010 2560 2030 2580
rect 2290 2560 2310 2580
rect 2570 2560 2590 2580
rect 2850 2560 2870 2580
rect 3130 2560 3150 2580
rect 3410 2560 3430 2580
rect 2010 2540 3430 2560
rect 1790 2520 1830 2530
rect 1930 2520 1970 2530
rect 3550 2520 3570 2580
rect 1790 2500 1800 2520
rect 1820 2500 1940 2520
rect 1960 2500 3570 2520
rect 1790 2490 1830 2500
rect 1930 2490 1970 2500
rect 2010 2460 3430 2480
rect 1790 2450 1830 2460
rect 1790 2430 1800 2450
rect 1820 2440 1830 2450
rect 2010 2440 2030 2460
rect 2290 2440 2310 2460
rect 2570 2440 2590 2460
rect 2850 2440 2870 2460
rect 3130 2440 3150 2460
rect 3410 2440 3430 2460
rect 3550 2440 3570 2500
rect 1820 2430 2040 2440
rect 1790 2420 2010 2430
rect 2000 2390 2010 2420
rect 2030 2390 2040 2430
rect 1790 2380 1830 2390
rect 2000 2380 2040 2390
rect 2140 2430 2180 2440
rect 2140 2390 2150 2430
rect 2170 2390 2180 2430
rect 2140 2380 2180 2390
rect 2280 2430 2320 2440
rect 2280 2390 2290 2430
rect 2310 2390 2320 2430
rect 2280 2380 2320 2390
rect 2420 2430 2460 2440
rect 2420 2390 2430 2430
rect 2450 2390 2460 2430
rect 2420 2380 2460 2390
rect 2560 2430 2600 2440
rect 2560 2390 2570 2430
rect 2590 2390 2600 2430
rect 2560 2380 2600 2390
rect 2700 2430 2740 2440
rect 2700 2390 2710 2430
rect 2730 2390 2740 2430
rect 2700 2380 2740 2390
rect 2840 2430 2880 2440
rect 2840 2390 2850 2430
rect 2870 2390 2880 2430
rect 2840 2380 2880 2390
rect 2980 2430 3020 2440
rect 2980 2390 2990 2430
rect 3010 2390 3020 2430
rect 2980 2380 3020 2390
rect 3120 2430 3160 2440
rect 3120 2390 3130 2430
rect 3150 2390 3160 2430
rect 3120 2380 3160 2390
rect 3260 2430 3300 2440
rect 3260 2390 3270 2430
rect 3290 2390 3300 2430
rect 3260 2380 3300 2390
rect 3400 2430 3440 2440
rect 3400 2390 3410 2430
rect 3430 2390 3440 2430
rect 3400 2380 3440 2390
rect 3540 2430 3620 2440
rect 3540 2390 3550 2430
rect 3570 2390 3590 2430
rect 3610 2390 3620 2430
rect 3540 2380 3620 2390
rect 1790 2360 1800 2380
rect 1820 2360 1830 2380
rect 1790 2350 1830 2360
rect 2150 2350 2170 2380
rect 2430 2350 2450 2380
rect 2710 2350 2730 2380
rect 2990 2350 3010 2380
rect 3270 2350 3290 2380
rect 1730 2340 1770 2350
rect 1730 2320 1740 2340
rect 1760 2320 1770 2340
rect 1730 2310 1770 2320
rect 1810 2340 1830 2350
rect 2140 2340 2180 2350
rect 2420 2340 2460 2350
rect 2700 2340 2740 2350
rect 2980 2340 3020 2350
rect 3260 2340 3300 2350
rect 1810 2320 2150 2340
rect 2170 2320 2430 2340
rect 2450 2320 2710 2340
rect 2730 2320 2990 2340
rect 3010 2320 3270 2340
rect 3290 2320 3300 2340
rect 1810 2290 1830 2320
rect 2140 2310 2180 2320
rect 2420 2310 2460 2320
rect 2700 2310 2740 2320
rect 2980 2310 3020 2320
rect 3260 2310 3300 2320
rect 3410 2320 3430 2380
rect 3550 2350 3570 2380
rect 3540 2340 3580 2350
rect 3540 2320 3550 2340
rect 3570 2320 3580 2340
rect 3410 2300 3510 2320
rect 3540 2310 3580 2320
rect 1770 2280 1830 2290
rect 1940 2280 2000 2290
rect 2110 2280 2170 2290
rect 2280 2280 2340 2290
rect 2450 2280 2510 2290
rect 2620 2280 2680 2290
rect 2790 2280 2850 2290
rect 2960 2280 3020 2290
rect 3130 2280 3190 2290
rect 3300 2280 3360 2290
rect 1770 2260 1780 2280
rect 1820 2260 1950 2280
rect 1990 2260 2120 2280
rect 2160 2260 2290 2280
rect 2330 2260 2460 2280
rect 2500 2260 2630 2280
rect 2670 2260 2800 2280
rect 2840 2260 2970 2280
rect 3010 2260 3140 2280
rect 3180 2260 3310 2280
rect 3350 2260 3460 2280
rect 1770 2250 1830 2260
rect 1940 2250 2000 2260
rect 2110 2250 2170 2260
rect 2280 2250 2340 2260
rect 2450 2250 2510 2260
rect 2620 2250 2680 2260
rect 2790 2250 2850 2260
rect 2960 2250 3020 2260
rect 3130 2250 3190 2260
rect 3300 2250 3360 2260
rect 3440 2180 3460 2260
rect 3430 2170 3470 2180
rect 3430 2150 3440 2170
rect 3460 2150 3470 2170
rect 3430 2140 3470 2150
rect 1770 2110 1830 2120
rect 1770 2090 1780 2110
rect 1820 2090 1830 2110
rect 1940 2110 2000 2120
rect 1940 2090 1950 2110
rect 1990 2090 2000 2110
rect 2110 2110 2170 2120
rect 2110 2090 2120 2110
rect 2160 2090 2170 2110
rect 2280 2110 2340 2120
rect 2280 2090 2290 2110
rect 2330 2090 2340 2110
rect 2450 2110 2510 2120
rect 2450 2090 2460 2110
rect 2500 2090 2510 2110
rect 2620 2110 2680 2120
rect 2620 2090 2630 2110
rect 2670 2090 2680 2110
rect 2790 2110 2850 2120
rect 2790 2090 2800 2110
rect 2840 2090 2850 2110
rect 2960 2110 3020 2120
rect 2960 2090 2970 2110
rect 3010 2090 3020 2110
rect 3130 2110 3190 2120
rect 3130 2090 3140 2110
rect 3180 2090 3190 2110
rect 3300 2110 3360 2120
rect 3300 2090 3310 2110
rect 3350 2090 3360 2110
rect 20 2070 3360 2090
rect 20 2050 30 2070
rect 70 2050 80 2070
rect 20 2040 80 2050
rect 190 2050 200 2070
rect 240 2050 250 2070
rect 190 2040 250 2050
rect 360 2050 370 2070
rect 410 2050 420 2070
rect 360 2040 420 2050
rect 530 2050 540 2070
rect 580 2050 590 2070
rect 530 2040 590 2050
rect 700 2050 710 2070
rect 750 2050 760 2070
rect 700 2040 760 2050
rect 870 2050 880 2070
rect 920 2050 930 2070
rect 870 2040 930 2050
rect 1040 2050 1050 2070
rect 1090 2050 1100 2070
rect 1040 2040 1100 2050
rect 1210 2050 1220 2070
rect 1260 2050 1270 2070
rect 1210 2040 1270 2050
rect 1380 2050 1390 2070
rect 1430 2050 1440 2070
rect 1380 2040 1440 2050
rect 1550 2050 1560 2070
rect 1600 2050 1610 2070
rect 1550 2040 1610 2050
rect -210 1550 -200 1570
rect -160 1550 -110 1570
rect -210 1540 -150 1550
rect -210 1030 -150 1040
rect -210 1010 -200 1030
rect -160 1010 -150 1030
rect -210 1000 -150 1010
rect 20 1030 80 1040
rect 20 1010 30 1030
rect 70 1010 80 1030
rect 20 1000 80 1010
rect 190 1030 250 1040
rect 190 1010 200 1030
rect 240 1010 250 1030
rect 190 1000 250 1010
rect 360 1030 420 1040
rect 360 1010 370 1030
rect 410 1010 420 1030
rect 360 1000 420 1010
rect 530 1030 590 1040
rect 530 1010 540 1030
rect 580 1010 590 1030
rect 530 1000 590 1010
rect 700 1030 760 1040
rect 700 1010 710 1030
rect 750 1010 760 1030
rect 700 1000 760 1010
rect 870 1030 930 1040
rect 870 1010 880 1030
rect 920 1010 930 1030
rect 870 1000 930 1010
rect 1040 1030 1100 1040
rect 1040 1010 1050 1030
rect 1090 1010 1100 1030
rect 1040 1000 1100 1010
rect 1210 1030 1270 1040
rect 1210 1010 1220 1030
rect 1260 1010 1270 1030
rect 1210 1000 1270 1010
rect 1380 1030 1440 1040
rect 1380 1010 1390 1030
rect 1430 1010 1440 1030
rect 1380 1000 1440 1010
rect 1550 1030 1610 1040
rect 1550 1010 1560 1030
rect 1600 1010 1610 1030
rect 1550 1000 1610 1010
rect -310 970 -270 980
rect -190 970 -170 1000
rect -310 950 -300 970
rect -280 950 -170 970
rect -310 940 -270 950
rect 20 -10 80 0
rect -60 -30 -20 -20
rect 20 -30 30 -10
rect 70 -30 80 -10
rect 190 -10 250 0
rect 190 -30 200 -10
rect 240 -30 250 -10
rect 360 -10 420 0
rect 360 -30 370 -10
rect 410 -30 420 -10
rect 530 -10 590 0
rect 530 -30 540 -10
rect 580 -30 590 -10
rect 700 -10 760 0
rect 700 -30 710 -10
rect 750 -30 760 -10
rect 870 -10 930 0
rect 870 -30 880 -10
rect 920 -30 930 -10
rect 1040 -10 1100 0
rect 1040 -30 1050 -10
rect 1090 -30 1100 -10
rect 1210 -10 1270 0
rect 1210 -30 1220 -10
rect 1260 -30 1270 -10
rect 1380 -10 1440 0
rect 1380 -30 1390 -10
rect 1430 -30 1440 -10
rect 1550 -10 1610 0
rect 1550 -30 1560 -10
rect 1600 -30 1610 -10
rect 1680 -30 1700 2070
rect 1770 2050 1780 2070
rect 1820 2050 1830 2070
rect 1770 2040 1830 2050
rect 1940 2050 1950 2070
rect 1990 2050 2000 2070
rect 1940 2040 2000 2050
rect 2110 2050 2120 2070
rect 2160 2050 2170 2070
rect 2110 2040 2170 2050
rect 2280 2050 2290 2070
rect 2330 2050 2340 2070
rect 2280 2040 2340 2050
rect 2450 2050 2460 2070
rect 2500 2050 2510 2070
rect 2450 2040 2510 2050
rect 2620 2050 2630 2070
rect 2670 2050 2680 2070
rect 2620 2040 2680 2050
rect 2790 2050 2800 2070
rect 2840 2050 2850 2070
rect 2790 2040 2850 2050
rect 2960 2050 2970 2070
rect 3010 2050 3020 2070
rect 2960 2040 3020 2050
rect 3130 2050 3140 2070
rect 3180 2050 3190 2070
rect 3130 2040 3190 2050
rect 3300 2050 3310 2070
rect 3350 2050 3360 2070
rect 3300 2040 3360 2050
rect 3490 1570 3510 2300
rect 3550 2120 3570 2310
rect 3530 2110 3590 2120
rect 3530 2090 3540 2110
rect 3580 2090 3590 2110
rect 3530 2080 3590 2090
rect 3530 1570 3590 1580
rect 3490 1550 3540 1570
rect 3580 1550 3590 1570
rect 3530 1540 3590 1550
rect 1770 1030 1830 1040
rect 1770 1010 1780 1030
rect 1820 1010 1830 1030
rect 1770 1000 1830 1010
rect 1940 1030 2000 1040
rect 1940 1010 1950 1030
rect 1990 1010 2000 1030
rect 1940 1000 2000 1010
rect 2110 1030 2170 1040
rect 2110 1010 2120 1030
rect 2160 1010 2170 1030
rect 2110 1000 2170 1010
rect 2280 1030 2340 1040
rect 2280 1010 2290 1030
rect 2330 1010 2340 1030
rect 2280 1000 2340 1010
rect 2450 1030 2510 1040
rect 2450 1010 2460 1030
rect 2500 1010 2510 1030
rect 2450 1000 2510 1010
rect 2620 1030 2680 1040
rect 2620 1010 2630 1030
rect 2670 1010 2680 1030
rect 2620 1000 2680 1010
rect 2790 1030 2850 1040
rect 2790 1010 2800 1030
rect 2840 1010 2850 1030
rect 2790 1000 2850 1010
rect 2960 1030 3020 1040
rect 2960 1010 2970 1030
rect 3010 1010 3020 1030
rect 2960 1000 3020 1010
rect 3130 1030 3190 1040
rect 3130 1010 3140 1030
rect 3180 1010 3190 1030
rect 3130 1000 3190 1010
rect 3300 1030 3360 1040
rect 3300 1010 3310 1030
rect 3350 1010 3360 1030
rect 3300 1000 3360 1010
rect 3530 1030 3590 1040
rect 3530 1010 3540 1030
rect 3580 1010 3590 1030
rect 3530 1000 3590 1010
rect 3550 970 3570 1000
rect 3660 980 3680 4040
rect 3650 970 3690 980
rect 3550 950 3660 970
rect 3680 950 3690 970
rect 3650 940 3690 950
rect 1770 -10 1830 0
rect 1770 -30 1780 -10
rect 1820 -30 1830 -10
rect 1940 -10 2000 0
rect 1940 -30 1950 -10
rect 1990 -30 2000 -10
rect 2110 -10 2170 0
rect 2110 -30 2120 -10
rect 2160 -30 2170 -10
rect 2280 -10 2340 0
rect 2280 -30 2290 -10
rect 2330 -30 2340 -10
rect 2450 -10 2510 0
rect 2450 -30 2460 -10
rect 2500 -30 2510 -10
rect 2620 -10 2680 0
rect 2620 -30 2630 -10
rect 2670 -30 2680 -10
rect 2790 -10 2850 0
rect 2790 -30 2800 -10
rect 2840 -30 2850 -10
rect 2960 -10 3020 0
rect 2960 -30 2970 -10
rect 3010 -30 3020 -10
rect 3130 -10 3190 0
rect 3130 -30 3140 -10
rect 3180 -30 3190 -10
rect 3300 -10 3360 0
rect 3300 -30 3310 -10
rect 3350 -30 3360 -10
rect 3400 -30 3440 -20
rect -60 -50 -50 -30
rect -30 -50 3410 -30
rect 3430 -50 3440 -30
rect -60 -60 -20 -50
rect 20 -70 30 -50
rect 70 -70 80 -50
rect 190 -70 200 -50
rect 240 -70 250 -50
rect 360 -70 370 -50
rect 410 -70 420 -50
rect 530 -70 540 -50
rect 580 -70 590 -50
rect 700 -70 710 -50
rect 750 -70 760 -50
rect 870 -70 880 -50
rect 920 -70 930 -50
rect 1040 -70 1050 -50
rect 1090 -70 1100 -50
rect 1210 -70 1220 -50
rect 1260 -70 1270 -50
rect 1380 -70 1390 -50
rect 1430 -70 1440 -50
rect 1550 -70 1560 -50
rect 1600 -70 1610 -50
rect 1770 -70 1780 -50
rect 1820 -70 1830 -50
rect 1940 -70 1950 -50
rect 1990 -70 2000 -50
rect 2110 -70 2120 -50
rect 2160 -70 2170 -50
rect 2280 -70 2290 -50
rect 2330 -70 2340 -50
rect 2450 -70 2460 -50
rect 2500 -70 2510 -50
rect 2620 -70 2630 -50
rect 2670 -70 2680 -50
rect 2790 -70 2800 -50
rect 2840 -70 2850 -50
rect 2960 -70 2970 -50
rect 3010 -70 3020 -50
rect 3130 -70 3140 -50
rect 3180 -70 3190 -50
rect 3300 -70 3310 -50
rect 3350 -70 3360 -50
rect 3400 -60 3440 -50
<< end >>
