magic
tech sky130A
timestamp 1762117721
<< nwell >>
rect -220 -460 300 170
rect 1280 -460 1800 170
<< nmos >>
rect 385 0 485 100
rect 615 0 715 100
rect 865 0 965 100
rect 1095 0 1195 100
rect 385 -130 485 -30
rect 615 -130 715 -30
rect 865 -130 965 -30
rect 1095 -130 1195 -30
rect 385 -260 485 -160
rect 615 -260 715 -160
rect 865 -260 965 -160
rect 1095 -260 1195 -160
rect 385 -390 485 -290
rect 615 -390 715 -290
rect 865 -390 965 -290
rect 1095 -390 1195 -290
<< pmos >>
rect -100 0 0 100
rect 130 0 230 100
rect 1350 0 1450 100
rect 1580 0 1680 100
rect -100 -130 0 -30
rect 130 -130 230 -30
rect 1350 -130 1450 -30
rect 1580 -130 1680 -30
rect -100 -260 0 -160
rect 130 -260 230 -160
rect 1350 -260 1450 -160
rect 1580 -260 1680 -160
rect -100 -390 0 -290
rect 130 -390 230 -290
rect 1350 -390 1450 -290
rect 1580 -390 1680 -290
<< ndiff >>
rect 335 85 385 100
rect 335 15 350 85
rect 370 15 385 85
rect 335 0 385 15
rect 485 85 535 100
rect 485 15 500 85
rect 520 15 535 85
rect 485 0 535 15
rect 565 85 615 100
rect 565 15 580 85
rect 600 15 615 85
rect 565 0 615 15
rect 715 85 765 100
rect 715 15 730 85
rect 750 15 765 85
rect 715 0 765 15
rect 815 85 865 100
rect 815 15 830 85
rect 850 15 865 85
rect 815 0 865 15
rect 965 85 1015 100
rect 965 15 980 85
rect 1000 15 1015 85
rect 965 0 1015 15
rect 1045 85 1095 100
rect 1045 15 1060 85
rect 1080 15 1095 85
rect 1045 0 1095 15
rect 1195 85 1245 100
rect 1195 15 1210 85
rect 1230 15 1245 85
rect 1195 0 1245 15
rect 335 -45 385 -30
rect 335 -115 350 -45
rect 370 -115 385 -45
rect 335 -130 385 -115
rect 485 -45 535 -30
rect 485 -115 500 -45
rect 520 -115 535 -45
rect 485 -130 535 -115
rect 565 -45 615 -30
rect 565 -115 580 -45
rect 600 -115 615 -45
rect 565 -130 615 -115
rect 715 -45 765 -30
rect 715 -115 730 -45
rect 750 -115 765 -45
rect 715 -130 765 -115
rect 815 -45 865 -30
rect 815 -115 830 -45
rect 850 -115 865 -45
rect 815 -130 865 -115
rect 965 -45 1015 -30
rect 965 -115 980 -45
rect 1000 -115 1015 -45
rect 965 -130 1015 -115
rect 1045 -45 1095 -30
rect 1045 -115 1060 -45
rect 1080 -115 1095 -45
rect 1045 -130 1095 -115
rect 1195 -45 1245 -30
rect 1195 -115 1210 -45
rect 1230 -115 1245 -45
rect 1195 -130 1245 -115
rect 335 -175 385 -160
rect 335 -245 350 -175
rect 370 -245 385 -175
rect 335 -260 385 -245
rect 485 -175 535 -160
rect 485 -245 500 -175
rect 520 -245 535 -175
rect 485 -260 535 -245
rect 565 -175 615 -160
rect 565 -245 580 -175
rect 600 -245 615 -175
rect 565 -260 615 -245
rect 715 -175 765 -160
rect 715 -245 730 -175
rect 750 -245 765 -175
rect 715 -260 765 -245
rect 815 -175 865 -160
rect 815 -245 830 -175
rect 850 -245 865 -175
rect 815 -260 865 -245
rect 965 -175 1015 -160
rect 965 -245 980 -175
rect 1000 -245 1015 -175
rect 965 -260 1015 -245
rect 1045 -175 1095 -160
rect 1045 -245 1060 -175
rect 1080 -245 1095 -175
rect 1045 -260 1095 -245
rect 1195 -175 1245 -160
rect 1195 -245 1210 -175
rect 1230 -245 1245 -175
rect 1195 -260 1245 -245
rect 335 -305 385 -290
rect 335 -375 350 -305
rect 370 -375 385 -305
rect 335 -390 385 -375
rect 485 -305 535 -290
rect 485 -375 500 -305
rect 520 -375 535 -305
rect 485 -390 535 -375
rect 565 -305 615 -290
rect 565 -375 580 -305
rect 600 -375 615 -305
rect 565 -390 615 -375
rect 715 -305 765 -290
rect 815 -305 865 -290
rect 715 -375 730 -305
rect 750 -375 765 -305
rect 815 -375 830 -305
rect 850 -375 865 -305
rect 715 -390 765 -375
rect 815 -390 865 -375
rect 965 -305 1015 -290
rect 965 -375 980 -305
rect 1000 -375 1015 -305
rect 965 -390 1015 -375
rect 1045 -305 1095 -290
rect 1045 -375 1060 -305
rect 1080 -375 1095 -305
rect 1045 -390 1095 -375
rect 1195 -305 1245 -290
rect 1195 -375 1210 -305
rect 1230 -375 1245 -305
rect 1195 -390 1245 -375
<< pdiff >>
rect -150 85 -100 100
rect -150 15 -135 85
rect -115 15 -100 85
rect -150 0 -100 15
rect 0 85 50 100
rect 0 15 15 85
rect 35 15 50 85
rect 0 0 50 15
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
rect 230 85 280 100
rect 230 15 245 85
rect 265 15 280 85
rect 230 0 280 15
rect 1300 85 1350 100
rect 1300 15 1315 85
rect 1335 15 1350 85
rect 1300 0 1350 15
rect 1450 85 1500 100
rect 1450 15 1465 85
rect 1485 15 1500 85
rect 1450 0 1500 15
rect 1530 85 1580 100
rect 1530 15 1545 85
rect 1565 15 1580 85
rect 1530 0 1580 15
rect 1680 85 1730 100
rect 1680 15 1695 85
rect 1715 15 1730 85
rect 1680 0 1730 15
rect -150 -45 -100 -30
rect -150 -115 -135 -45
rect -115 -115 -100 -45
rect -150 -130 -100 -115
rect 0 -45 50 -30
rect 0 -115 15 -45
rect 35 -115 50 -45
rect 0 -130 50 -115
rect 80 -45 130 -30
rect 80 -115 95 -45
rect 115 -115 130 -45
rect 80 -130 130 -115
rect 230 -45 280 -30
rect 230 -115 245 -45
rect 265 -115 280 -45
rect 230 -130 280 -115
rect 1300 -45 1350 -30
rect 1300 -115 1315 -45
rect 1335 -115 1350 -45
rect 1300 -130 1350 -115
rect 1450 -45 1500 -30
rect 1450 -115 1465 -45
rect 1485 -115 1500 -45
rect 1450 -130 1500 -115
rect 1530 -45 1580 -30
rect 1530 -115 1545 -45
rect 1565 -115 1580 -45
rect 1530 -130 1580 -115
rect 1680 -45 1730 -30
rect 1680 -115 1695 -45
rect 1715 -115 1730 -45
rect 1680 -130 1730 -115
rect -150 -175 -100 -160
rect -150 -245 -135 -175
rect -115 -245 -100 -175
rect -150 -260 -100 -245
rect 0 -175 50 -160
rect 0 -245 15 -175
rect 35 -245 50 -175
rect 0 -260 50 -245
rect 80 -175 130 -160
rect 80 -245 95 -175
rect 115 -245 130 -175
rect 80 -260 130 -245
rect 230 -175 280 -160
rect 230 -245 245 -175
rect 265 -245 280 -175
rect 230 -260 280 -245
rect 1300 -175 1350 -160
rect 1300 -245 1315 -175
rect 1335 -245 1350 -175
rect 1300 -260 1350 -245
rect 1450 -175 1500 -160
rect 1450 -245 1465 -175
rect 1485 -245 1500 -175
rect 1450 -260 1500 -245
rect 1530 -175 1580 -160
rect 1530 -245 1545 -175
rect 1565 -245 1580 -175
rect 1530 -260 1580 -245
rect 1680 -175 1730 -160
rect 1680 -245 1695 -175
rect 1715 -245 1730 -175
rect 1680 -260 1730 -245
rect -150 -305 -100 -290
rect -150 -375 -135 -305
rect -115 -375 -100 -305
rect -150 -390 -100 -375
rect 0 -305 50 -290
rect 0 -375 15 -305
rect 35 -375 50 -305
rect 0 -390 50 -375
rect 80 -305 130 -290
rect 80 -375 95 -305
rect 115 -375 130 -305
rect 80 -390 130 -375
rect 230 -305 280 -290
rect 230 -375 245 -305
rect 265 -375 280 -305
rect 230 -390 280 -375
rect 1300 -305 1350 -290
rect 1300 -375 1315 -305
rect 1335 -375 1350 -305
rect 1300 -390 1350 -375
rect 1450 -305 1500 -290
rect 1450 -375 1465 -305
rect 1485 -375 1500 -305
rect 1450 -390 1500 -375
rect 1530 -305 1580 -290
rect 1530 -375 1545 -305
rect 1565 -375 1580 -305
rect 1530 -390 1580 -375
rect 1680 -305 1730 -290
rect 1680 -375 1695 -305
rect 1715 -375 1730 -305
rect 1680 -390 1730 -375
<< ndiffc >>
rect 350 15 370 85
rect 500 15 520 85
rect 580 15 600 85
rect 730 15 750 85
rect 830 15 850 85
rect 980 15 1000 85
rect 1060 15 1080 85
rect 1210 15 1230 85
rect 350 -115 370 -45
rect 500 -115 520 -45
rect 580 -115 600 -45
rect 730 -115 750 -45
rect 830 -115 850 -45
rect 980 -115 1000 -45
rect 1060 -115 1080 -45
rect 1210 -115 1230 -45
rect 350 -245 370 -175
rect 500 -245 520 -175
rect 580 -245 600 -175
rect 730 -245 750 -175
rect 830 -245 850 -175
rect 980 -245 1000 -175
rect 1060 -245 1080 -175
rect 1210 -245 1230 -175
rect 350 -375 370 -305
rect 500 -375 520 -305
rect 580 -375 600 -305
rect 730 -375 750 -305
rect 830 -375 850 -305
rect 980 -375 1000 -305
rect 1060 -375 1080 -305
rect 1210 -375 1230 -305
<< pdiffc >>
rect -135 15 -115 85
rect 15 15 35 85
rect 95 15 115 85
rect 245 15 265 85
rect 1315 15 1335 85
rect 1465 15 1485 85
rect 1545 15 1565 85
rect 1695 15 1715 85
rect -135 -115 -115 -45
rect 15 -115 35 -45
rect 95 -115 115 -45
rect 245 -115 265 -45
rect 1315 -115 1335 -45
rect 1465 -115 1485 -45
rect 1545 -115 1565 -45
rect 1695 -115 1715 -45
rect -135 -245 -115 -175
rect 15 -245 35 -175
rect 95 -245 115 -175
rect 245 -245 265 -175
rect 1315 -245 1335 -175
rect 1465 -245 1485 -175
rect 1545 -245 1565 -175
rect 1695 -245 1715 -175
rect -135 -375 -115 -305
rect 15 -375 35 -305
rect 95 -375 115 -305
rect 245 -375 265 -305
rect 1315 -375 1335 -305
rect 1465 -375 1485 -305
rect 1545 -375 1565 -305
rect 1695 -375 1715 -305
<< psubdiff >>
rect 765 -305 815 -290
rect 765 -375 780 -305
rect 800 -375 815 -305
rect 765 -390 815 -375
<< nsubdiff >>
rect -200 85 -150 100
rect -200 15 -185 85
rect -165 15 -150 85
rect -200 0 -150 15
rect 1730 85 1780 100
rect 1730 15 1745 85
rect 1765 15 1780 85
rect 1730 0 1780 15
<< psubdiffcont >>
rect 780 -375 800 -305
<< nsubdiffcont >>
rect -185 15 -165 85
rect 1745 15 1765 85
<< poly >>
rect 130 160 170 170
rect 130 140 140 160
rect 160 140 170 160
rect 130 130 170 140
rect 615 160 655 170
rect 615 140 625 160
rect 645 140 655 160
rect 615 130 655 140
rect 925 160 965 170
rect 925 140 935 160
rect 955 140 965 160
rect 925 130 965 140
rect 1410 160 1450 170
rect 1410 140 1420 160
rect 1440 140 1450 160
rect 1410 130 1450 140
rect -100 100 0 130
rect 130 100 230 130
rect 385 100 485 130
rect 615 100 715 130
rect 865 100 965 130
rect 1095 100 1195 130
rect 1350 100 1450 130
rect 1580 100 1680 130
rect -100 -30 0 0
rect 130 -30 230 0
rect 385 -30 485 0
rect 615 -30 715 0
rect 865 -30 965 0
rect 1095 -30 1195 0
rect 1350 -30 1450 0
rect 1580 -30 1680 0
rect -100 -160 0 -130
rect 130 -160 230 -130
rect 385 -160 485 -130
rect 615 -160 715 -130
rect 865 -160 965 -130
rect 1095 -160 1195 -130
rect 1350 -160 1450 -130
rect 1580 -160 1680 -130
rect -100 -290 0 -260
rect 130 -290 230 -260
rect 385 -290 485 -260
rect 615 -290 715 -260
rect 865 -290 965 -260
rect 1095 -290 1195 -260
rect 1350 -290 1450 -260
rect 1580 -290 1680 -260
rect -100 -420 0 -390
rect 130 -420 230 -390
rect -40 -430 0 -420
rect -40 -450 -30 -430
rect -10 -450 0 -430
rect -40 -460 0 -450
rect 190 -430 230 -420
rect 190 -450 200 -430
rect 220 -450 230 -430
rect 190 -460 230 -450
rect 385 -420 485 -390
rect 615 -420 715 -390
rect 385 -430 425 -420
rect 385 -450 395 -430
rect 415 -450 425 -430
rect 385 -460 425 -450
rect 675 -430 715 -420
rect 675 -450 685 -430
rect 705 -450 715 -430
rect 675 -460 715 -450
rect 865 -420 965 -390
rect 1095 -420 1195 -390
rect 865 -430 905 -420
rect 865 -450 875 -430
rect 895 -450 905 -430
rect 865 -460 905 -450
rect 1155 -430 1195 -420
rect 1155 -450 1165 -430
rect 1185 -450 1195 -430
rect 1155 -460 1195 -450
rect 1350 -420 1450 -390
rect 1580 -420 1680 -390
rect 1350 -430 1390 -420
rect 1350 -450 1360 -430
rect 1380 -450 1390 -430
rect 1350 -460 1390 -450
rect 1580 -430 1620 -420
rect 1580 -450 1590 -430
rect 1610 -450 1620 -430
rect 1580 -460 1620 -450
<< polycont >>
rect 140 140 160 160
rect 625 140 645 160
rect 935 140 955 160
rect 1420 140 1440 160
rect -30 -450 -10 -430
rect 200 -450 220 -430
rect 395 -450 415 -430
rect 685 -450 705 -430
rect 875 -450 895 -430
rect 1165 -450 1185 -430
rect 1360 -450 1380 -430
rect 1590 -450 1610 -430
<< locali >>
rect 130 190 1820 210
rect 130 170 170 190
rect 1410 170 1450 190
rect 5 160 170 170
rect 5 140 140 160
rect 160 140 170 160
rect 5 130 170 140
rect 235 160 655 170
rect 235 140 625 160
rect 645 140 655 160
rect 235 130 655 140
rect 925 160 1345 170
rect 925 140 935 160
rect 955 140 1345 160
rect 925 130 1345 140
rect 1410 160 1575 170
rect 1410 140 1420 160
rect 1440 140 1575 160
rect 1410 130 1575 140
rect -195 85 -105 95
rect -195 15 -185 85
rect -165 15 -135 85
rect -115 15 -105 85
rect -195 5 -105 15
rect -145 -45 -105 5
rect -145 -115 -135 -45
rect -115 -115 -105 -45
rect -145 -175 -105 -115
rect 5 85 45 130
rect 5 15 15 85
rect 35 15 45 85
rect 5 -45 45 15
rect 5 -115 15 -45
rect 35 -115 45 -45
rect 5 -125 45 -115
rect 85 85 125 95
rect 85 15 95 85
rect 115 15 125 85
rect 85 -45 125 15
rect 85 -115 95 -45
rect 115 -115 125 -45
rect -145 -245 -135 -175
rect -115 -245 -105 -175
rect -145 -305 -105 -245
rect -145 -375 -135 -305
rect -115 -375 -105 -305
rect -145 -385 -105 -375
rect 5 -175 45 -165
rect 5 -245 15 -175
rect 35 -245 45 -175
rect 5 -305 45 -245
rect 5 -375 15 -305
rect 35 -375 45 -305
rect 5 -420 45 -375
rect 85 -175 125 -115
rect 235 85 275 130
rect 235 15 245 85
rect 265 15 275 85
rect 235 -45 275 15
rect 235 -115 245 -45
rect 265 -115 275 -45
rect 235 -125 275 -115
rect 340 85 380 95
rect 340 15 350 85
rect 370 15 380 85
rect 340 -45 380 15
rect 340 -115 350 -45
rect 370 -115 380 -45
rect 340 -125 380 -115
rect 490 85 530 95
rect 490 15 500 85
rect 520 15 530 85
rect 490 -45 530 15
rect 490 -115 500 -45
rect 520 -115 530 -45
rect 490 -125 530 -115
rect 570 85 610 130
rect 570 15 580 85
rect 600 15 610 85
rect 570 -45 610 15
rect 570 -115 580 -45
rect 600 -115 610 -45
rect 570 -125 610 -115
rect 720 85 760 95
rect 720 15 730 85
rect 750 15 760 85
rect 720 -45 760 15
rect 720 -115 730 -45
rect 750 -115 760 -45
rect 85 -245 95 -175
rect 115 -245 125 -175
rect 85 -305 125 -245
rect 85 -375 95 -305
rect 115 -375 125 -305
rect 85 -385 125 -375
rect 235 -175 275 -165
rect 235 -245 245 -175
rect 265 -245 275 -175
rect 235 -260 275 -245
rect 340 -175 380 -165
rect 340 -245 350 -175
rect 370 -245 380 -175
rect 340 -260 380 -245
rect 235 -290 380 -260
rect 235 -305 275 -290
rect 235 -375 245 -305
rect 265 -375 275 -305
rect 235 -385 275 -375
rect 340 -305 380 -290
rect 340 -375 350 -305
rect 370 -375 380 -305
rect 340 -420 380 -375
rect 490 -175 530 -165
rect 490 -245 500 -175
rect 520 -245 530 -175
rect 490 -305 530 -245
rect 490 -375 500 -305
rect 520 -375 530 -305
rect 490 -390 530 -375
rect 570 -175 610 -160
rect 570 -245 580 -175
rect 600 -245 610 -175
rect 570 -305 610 -245
rect 570 -375 580 -305
rect 600 -375 610 -305
rect -40 -430 45 -420
rect -40 -450 -30 -430
rect -10 -450 45 -430
rect -40 -460 45 -450
rect 190 -430 230 -420
rect 190 -450 200 -430
rect 220 -450 230 -430
rect 190 -480 230 -450
rect 340 -430 425 -420
rect 340 -450 395 -430
rect 415 -450 425 -430
rect 340 -460 425 -450
rect 570 -480 610 -375
rect 720 -175 760 -115
rect 720 -245 730 -175
rect 750 -245 760 -175
rect 720 -295 760 -245
rect 820 85 860 95
rect 820 15 830 85
rect 850 15 860 85
rect 820 -45 860 15
rect 820 -115 830 -45
rect 850 -115 860 -45
rect 820 -175 860 -115
rect 970 85 1010 130
rect 970 15 980 85
rect 1000 15 1010 85
rect 970 -45 1010 15
rect 970 -115 980 -45
rect 1000 -115 1010 -45
rect 970 -125 1010 -115
rect 1050 85 1090 95
rect 1050 15 1060 85
rect 1080 15 1090 85
rect 1050 -45 1090 15
rect 1050 -115 1060 -45
rect 1080 -115 1090 -45
rect 1050 -125 1090 -115
rect 1200 85 1240 95
rect 1200 15 1210 85
rect 1230 15 1240 85
rect 1200 -45 1240 15
rect 1200 -115 1210 -45
rect 1230 -115 1240 -45
rect 1200 -125 1240 -115
rect 1305 85 1345 130
rect 1305 15 1315 85
rect 1335 15 1345 85
rect 1305 -45 1345 15
rect 1305 -115 1315 -45
rect 1335 -115 1345 -45
rect 1305 -125 1345 -115
rect 1455 85 1495 95
rect 1455 15 1465 85
rect 1485 15 1495 85
rect 1455 -45 1495 15
rect 1455 -115 1465 -45
rect 1485 -115 1495 -45
rect 820 -245 830 -175
rect 850 -245 860 -175
rect 820 -295 860 -245
rect 720 -305 860 -295
rect 720 -375 730 -305
rect 750 -375 780 -305
rect 800 -375 830 -305
rect 850 -375 860 -305
rect 720 -385 860 -375
rect 970 -175 1010 -160
rect 970 -245 980 -175
rect 1000 -245 1010 -175
rect 970 -305 1010 -245
rect 970 -375 980 -305
rect 1000 -375 1010 -305
rect 675 -430 905 -420
rect 675 -450 685 -430
rect 705 -450 875 -430
rect 895 -450 905 -430
rect 675 -460 905 -450
rect 190 -500 610 -480
rect 765 -520 815 -460
rect 970 -480 1010 -375
rect 1050 -175 1090 -165
rect 1050 -245 1060 -175
rect 1080 -245 1090 -175
rect 1050 -305 1090 -245
rect 1050 -375 1060 -305
rect 1080 -375 1090 -305
rect 1050 -390 1090 -375
rect 1200 -175 1240 -165
rect 1200 -245 1210 -175
rect 1230 -245 1240 -175
rect 1200 -260 1240 -245
rect 1305 -175 1345 -165
rect 1305 -245 1315 -175
rect 1335 -245 1345 -175
rect 1305 -260 1345 -245
rect 1200 -290 1345 -260
rect 1200 -305 1240 -290
rect 1200 -375 1210 -305
rect 1230 -375 1240 -305
rect 1200 -420 1240 -375
rect 1305 -305 1345 -290
rect 1305 -375 1315 -305
rect 1335 -375 1345 -305
rect 1305 -385 1345 -375
rect 1455 -175 1495 -115
rect 1535 85 1575 130
rect 1535 15 1545 85
rect 1565 15 1575 85
rect 1535 -45 1575 15
rect 1535 -115 1545 -45
rect 1565 -115 1575 -45
rect 1535 -125 1575 -115
rect 1685 85 1775 95
rect 1685 15 1695 85
rect 1715 15 1745 85
rect 1765 15 1775 85
rect 1685 5 1775 15
rect 1685 -45 1725 5
rect 1685 -115 1695 -45
rect 1715 -115 1725 -45
rect 1455 -245 1465 -175
rect 1485 -245 1495 -175
rect 1455 -305 1495 -245
rect 1455 -375 1465 -305
rect 1485 -375 1495 -305
rect 1455 -385 1495 -375
rect 1535 -175 1575 -165
rect 1535 -245 1545 -175
rect 1565 -245 1575 -175
rect 1535 -305 1575 -245
rect 1535 -375 1545 -305
rect 1565 -375 1575 -305
rect 1535 -420 1575 -375
rect 1685 -175 1725 -115
rect 1685 -245 1695 -175
rect 1715 -245 1725 -175
rect 1685 -305 1725 -245
rect 1685 -375 1695 -305
rect 1715 -375 1725 -305
rect 1685 -385 1725 -375
rect 1155 -430 1240 -420
rect 1155 -450 1165 -430
rect 1185 -450 1240 -430
rect 1155 -460 1240 -450
rect 1350 -430 1390 -420
rect 1350 -450 1360 -430
rect 1380 -450 1390 -430
rect 1350 -480 1390 -450
rect 1535 -430 1620 -420
rect 1535 -450 1590 -430
rect 1610 -450 1620 -430
rect 1535 -460 1620 -450
rect 970 -500 1390 -480
rect 765 -540 1820 -520
<< viali >>
rect -135 15 -115 85
rect 95 15 115 85
rect 15 -245 35 -175
rect 350 15 370 85
rect 350 -115 370 -45
rect 500 15 520 85
rect 730 15 750 85
rect 350 -245 370 -175
rect 500 -375 520 -305
rect 830 15 850 85
rect 1060 15 1080 85
rect 1210 15 1230 85
rect 1210 -115 1230 -45
rect 1465 15 1485 85
rect 780 -375 800 -305
rect 1060 -375 1080 -305
rect 1210 -245 1230 -175
rect 1695 15 1715 85
rect 1545 -245 1565 -175
<< metal1 >>
rect 85 130 1500 170
rect 85 95 125 130
rect -220 85 125 95
rect -220 15 -135 85
rect -115 15 95 85
rect 115 15 125 85
rect -220 0 125 15
rect 325 85 380 100
rect 325 15 340 85
rect 370 15 380 85
rect 325 0 380 15
rect 490 85 760 95
rect 490 15 500 85
rect 520 15 730 85
rect 750 15 760 85
rect 490 0 760 15
rect 820 85 1090 95
rect 820 15 830 85
rect 850 15 1060 85
rect 1080 15 1090 85
rect 820 0 1090 15
rect 1200 85 1245 100
rect 1200 15 1210 85
rect 1240 15 1245 85
rect 1200 0 1245 15
rect 1455 95 1500 130
rect 1455 85 1820 95
rect 1455 15 1465 85
rect 1485 15 1695 85
rect 1715 15 1820 85
rect 1455 0 1820 15
rect 5 -45 380 -30
rect 5 -115 350 -45
rect 370 -115 380 -45
rect 5 -130 380 -115
rect 1200 -45 1575 -30
rect 1200 -115 1210 -45
rect 1230 -115 1575 -45
rect 1200 -130 1575 -115
rect 5 -175 50 -130
rect 5 -245 15 -175
rect 35 -245 50 -175
rect 5 -260 50 -245
rect 335 -175 1245 -160
rect 335 -245 350 -175
rect 370 -245 1210 -175
rect 1230 -245 1245 -175
rect 335 -260 1245 -245
rect 1530 -175 1575 -130
rect 1530 -245 1545 -175
rect 1565 -245 1575 -175
rect 1530 -260 1575 -245
rect 490 -305 535 -290
rect 490 -375 500 -305
rect 530 -375 535 -305
rect 490 -560 535 -375
rect 765 -305 815 -295
rect 765 -375 780 -305
rect 800 -375 815 -305
rect 765 -540 815 -375
rect 1035 -305 1090 -290
rect 1035 -375 1050 -305
rect 1080 -375 1090 -305
rect 1035 -390 1090 -375
rect 765 -560 1820 -540
<< via1 >>
rect 340 15 350 85
rect 350 15 370 85
rect 1210 15 1230 85
rect 1230 15 1240 85
rect 500 -375 520 -305
rect 520 -375 530 -305
rect 1050 -375 1060 -305
rect 1060 -375 1080 -305
<< metal2 >>
rect 325 85 1245 100
rect 325 15 340 85
rect 370 15 1210 85
rect 1240 15 1245 85
rect 325 0 1245 15
rect 490 -305 1090 -290
rect 490 -375 500 -305
rect 530 -375 1050 -305
rect 1080 -375 1090 -305
rect 490 -390 1090 -375
<< labels >>
rlabel metal1 1820 50 1820 50 3 VP
port 1 e
rlabel locali 1820 200 1820 200 3 VBP
port 2 e
rlabel locali 1820 -530 1820 -530 3 VBN
port 3 e
rlabel metal1 1820 -550 1820 -550 3 VN
port 4 e
rlabel metal1 515 -560 515 -560 5 RES
port 5 s
<< end >>
