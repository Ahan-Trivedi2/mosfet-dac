magic
tech sky130A
timestamp 1762117972
<< nmos >>
rect -130 2755 -55 3255
rect 55 2755 130 3255
rect 410 2755 485 3255
rect 595 2755 670 3255
rect 950 2755 1025 3255
rect 1135 2755 1210 3255
rect 1490 2755 1565 3255
rect 1675 2755 1750 3255
rect 2030 2755 2105 3255
rect 2215 2755 2290 3255
rect 2570 2755 2645 3255
rect 2755 2755 2830 3255
rect 3110 2755 3185 3255
rect 3295 2755 3370 3255
rect -130 2205 -55 2705
rect 55 2205 130 2705
rect 410 2205 485 2705
rect 595 2205 670 2705
rect 950 2205 1025 2705
rect 1135 2205 1210 2705
rect 1490 2205 1565 2705
rect 1675 2205 1750 2705
rect 2030 2205 2105 2705
rect 2215 2205 2290 2705
rect 2570 2205 2645 2705
rect 2755 2205 2830 2705
rect 3110 2205 3185 2705
rect 3295 2205 3370 2705
rect -130 1655 -55 2155
rect 55 1655 130 2155
rect 410 1655 485 2155
rect 595 1655 670 2155
rect 950 1655 1025 2155
rect 1135 1655 1210 2155
rect 1490 1655 1565 2155
rect 1675 1655 1750 2155
rect 2030 1655 2105 2155
rect 2215 1655 2290 2155
rect 2570 1655 2645 2155
rect 2755 1655 2830 2155
rect 3110 1655 3185 2155
rect 3295 1655 3370 2155
rect -130 1105 -55 1605
rect 55 1105 130 1605
rect 410 1105 485 1605
rect 595 1105 670 1605
rect 950 1105 1025 1605
rect 1135 1105 1210 1605
rect 1490 1105 1565 1605
rect 1675 1105 1750 1605
rect 2030 1105 2105 1605
rect 2215 1105 2290 1605
rect 2570 1105 2645 1605
rect 2755 1105 2830 1605
rect 3110 1105 3185 1605
rect 3295 1105 3370 1605
rect -130 555 -55 1055
rect 55 555 130 1055
rect 410 555 485 1055
rect 595 555 670 1055
rect 950 555 1025 1055
rect 1135 555 1210 1055
rect 1490 555 1565 1055
rect 1675 555 1750 1055
rect 2030 555 2105 1055
rect 2215 555 2290 1055
rect 2570 555 2645 1055
rect 2755 555 2830 1055
rect 3110 555 3185 1055
rect 3295 555 3370 1055
rect -130 -125 -55 375
rect 55 -125 130 375
rect 410 -125 485 375
rect 595 -125 670 375
rect 950 -125 1025 375
rect 1135 -125 1210 375
rect 1490 -125 1565 375
rect 1675 -125 1750 375
rect 2030 -125 2105 375
rect 2215 -125 2290 375
rect 2570 -125 2645 375
rect 2755 -125 2830 375
rect 3110 -125 3185 375
rect 3295 -125 3370 375
rect 3650 -125 3725 375
rect -130 -675 -55 -175
rect 55 -675 130 -175
rect 410 -675 485 -175
rect 595 -675 670 -175
rect 950 -675 1025 -175
rect 1135 -675 1210 -175
rect 1490 -675 1565 -175
rect 1675 -675 1750 -175
rect 2030 -675 2105 -175
rect 2215 -675 2290 -175
rect 2570 -675 2645 -175
rect 2755 -675 2830 -175
rect 3110 -675 3185 -175
rect 3295 -675 3370 -175
rect 3650 -675 3725 -175
rect -130 -1225 -55 -725
rect 55 -1225 130 -725
rect 410 -1225 485 -725
rect 595 -1225 670 -725
rect 950 -1225 1025 -725
rect 1135 -1225 1210 -725
rect 1490 -1225 1565 -725
rect 1675 -1225 1750 -725
rect 2030 -1225 2105 -725
rect 2215 -1225 2290 -725
rect 2570 -1225 2645 -725
rect 2755 -1225 2830 -725
rect 3110 -1225 3185 -725
rect 3295 -1225 3370 -725
rect 3650 -1225 3725 -725
rect -130 -1775 -55 -1275
rect 55 -1775 130 -1275
rect 410 -1775 485 -1275
rect 595 -1775 670 -1275
rect 950 -1775 1025 -1275
rect 1135 -1775 1210 -1275
rect 1490 -1775 1565 -1275
rect 1675 -1775 1750 -1275
rect 2030 -1775 2105 -1275
rect 2215 -1775 2290 -1275
rect 2570 -1775 2645 -1275
rect 2755 -1775 2830 -1275
rect 3110 -1775 3185 -1275
rect 3295 -1775 3370 -1275
rect 3650 -1775 3725 -1275
rect -130 -2325 -55 -1825
rect 55 -2325 130 -1825
rect 410 -2325 485 -1825
rect 595 -2325 670 -1825
rect 950 -2325 1025 -1825
rect 1135 -2325 1210 -1825
rect 1490 -2325 1565 -1825
rect 1675 -2325 1750 -1825
rect 2030 -2325 2105 -1825
rect 2215 -2325 2290 -1825
rect 2570 -2325 2645 -1825
rect 2755 -2325 2830 -1825
rect 3110 -2325 3185 -1825
rect 3295 -2325 3370 -1825
rect 3650 -2325 3725 -1825
rect -130 -2960 -55 -2460
rect 55 -2960 130 -2460
rect 410 -2960 485 -2460
rect 595 -2960 670 -2460
rect 950 -2960 1025 -2460
rect 1135 -2960 1210 -2460
rect 1490 -2960 1565 -2460
rect 1675 -2960 1750 -2460
rect 2030 -2960 2105 -2460
rect 2215 -2960 2290 -2460
rect 2570 -2960 2645 -2460
rect 2755 -2960 2830 -2460
rect 3110 -2960 3185 -2460
rect 3295 -2960 3370 -2460
rect 3650 -2960 3725 -2460
rect -130 -3510 -55 -3010
rect 55 -3510 130 -3010
rect 410 -3510 485 -3010
rect 595 -3510 670 -3010
rect 950 -3510 1025 -3010
rect 1135 -3510 1210 -3010
rect 1490 -3510 1565 -3010
rect 1675 -3510 1750 -3010
rect 2030 -3510 2105 -3010
rect 2215 -3510 2290 -3010
rect 2570 -3510 2645 -3010
rect 2755 -3510 2830 -3010
rect 3110 -3510 3185 -3010
rect 3295 -3510 3370 -3010
rect 3650 -3510 3725 -3010
rect -130 -4060 -55 -3560
rect 55 -4060 130 -3560
rect 410 -4060 485 -3560
rect 595 -4060 670 -3560
rect 950 -4060 1025 -3560
rect 1135 -4060 1210 -3560
rect 1490 -4060 1565 -3560
rect 1675 -4060 1750 -3560
rect 2030 -4060 2105 -3560
rect 2215 -4060 2290 -3560
rect 2570 -4060 2645 -3560
rect 2755 -4060 2830 -3560
rect 3110 -4060 3185 -3560
rect 3295 -4060 3370 -3560
rect 3650 -4060 3725 -3560
rect -130 -4610 -55 -4110
rect 55 -4610 130 -4110
rect 410 -4610 485 -4110
rect 595 -4610 670 -4110
rect 950 -4610 1025 -4110
rect 1135 -4610 1210 -4110
rect 1490 -4610 1565 -4110
rect 1675 -4610 1750 -4110
rect 2030 -4610 2105 -4110
rect 2215 -4610 2290 -4110
rect 2570 -4610 2645 -4110
rect 2755 -4610 2830 -4110
rect 3110 -4610 3185 -4110
rect 3295 -4610 3370 -4110
rect 3650 -4610 3725 -4110
rect -130 -5160 -55 -4660
rect 55 -5160 130 -4660
rect 410 -5160 485 -4660
rect 595 -5160 670 -4660
rect 950 -5160 1025 -4660
rect 1135 -5160 1210 -4660
rect 1490 -5160 1565 -4660
rect 1675 -5160 1750 -4660
rect 2030 -5160 2105 -4660
rect 2215 -5160 2290 -4660
rect 2570 -5160 2645 -4660
rect 2755 -5160 2830 -4660
rect 3110 -5160 3185 -4660
rect 3295 -5160 3370 -4660
rect 3650 -5160 3725 -4660
rect -130 -5865 -55 -5365
rect 55 -5865 130 -5365
rect 410 -5865 485 -5365
rect 595 -5865 670 -5365
rect 950 -5865 1025 -5365
rect 1135 -5865 1210 -5365
rect 1490 -5865 1565 -5365
rect 1675 -5865 1750 -5365
rect 2030 -5865 2105 -5365
rect 2215 -5865 2290 -5365
rect 2570 -5865 2645 -5365
rect 2755 -5865 2830 -5365
rect 3110 -5865 3185 -5365
rect 3295 -5865 3370 -5365
rect -130 -6415 -55 -5915
rect 55 -6415 130 -5915
rect 410 -6415 485 -5915
rect 595 -6415 670 -5915
rect 950 -6415 1025 -5915
rect 1135 -6415 1210 -5915
rect 1490 -6415 1565 -5915
rect 1675 -6415 1750 -5915
rect 2030 -6415 2105 -5915
rect 2215 -6415 2290 -5915
rect 2570 -6415 2645 -5915
rect 2755 -6415 2830 -5915
rect 3110 -6415 3185 -5915
rect 3295 -6415 3370 -5915
rect -130 -6965 -55 -6465
rect 55 -6965 130 -6465
rect 410 -6965 485 -6465
rect 595 -6965 670 -6465
rect 950 -6965 1025 -6465
rect 1135 -6965 1210 -6465
rect 1490 -6965 1565 -6465
rect 1675 -6965 1750 -6465
rect 2030 -6965 2105 -6465
rect 2215 -6965 2290 -6465
rect 2570 -6965 2645 -6465
rect 2755 -6965 2830 -6465
rect 3110 -6965 3185 -6465
rect 3295 -6965 3370 -6465
rect -130 -7515 -55 -7015
rect 55 -7515 130 -7015
rect 410 -7515 485 -7015
rect 595 -7515 670 -7015
rect 950 -7515 1025 -7015
rect 1135 -7515 1210 -7015
rect 1490 -7515 1565 -7015
rect 1675 -7515 1750 -7015
rect 2030 -7515 2105 -7015
rect 2215 -7515 2290 -7015
rect 2570 -7515 2645 -7015
rect 2755 -7515 2830 -7015
rect 3110 -7515 3185 -7015
rect 3295 -7515 3370 -7015
rect -130 -8065 -55 -7565
rect 55 -8065 130 -7565
rect 410 -8065 485 -7565
rect 595 -8065 670 -7565
rect 950 -8065 1025 -7565
rect 1135 -8065 1210 -7565
rect 1490 -8065 1565 -7565
rect 1675 -8065 1750 -7565
rect 2030 -8065 2105 -7565
rect 2215 -8065 2290 -7565
rect 2570 -8065 2645 -7565
rect 2755 -8065 2830 -7565
rect 3110 -8065 3185 -7565
rect 3295 -8065 3370 -7565
<< ndiff >>
rect -130 3290 -55 3305
rect -130 3270 -115 3290
rect -70 3270 -55 3290
rect -130 3255 -55 3270
rect 55 3290 130 3305
rect 55 3270 70 3290
rect 115 3270 130 3290
rect 55 3255 130 3270
rect 410 3290 485 3305
rect 410 3270 425 3290
rect 470 3270 485 3290
rect 410 3255 485 3270
rect 595 3290 670 3305
rect 595 3270 610 3290
rect 655 3270 670 3290
rect 595 3255 670 3270
rect 950 3290 1025 3305
rect 950 3270 965 3290
rect 1010 3270 1025 3290
rect 950 3255 1025 3270
rect 1135 3290 1210 3305
rect 1135 3270 1150 3290
rect 1195 3270 1210 3290
rect 1135 3255 1210 3270
rect 1490 3290 1565 3305
rect 1490 3270 1505 3290
rect 1550 3270 1565 3290
rect 1490 3255 1565 3270
rect 1675 3290 1750 3305
rect 1675 3270 1690 3290
rect 1735 3270 1750 3290
rect 1675 3255 1750 3270
rect 2030 3290 2105 3305
rect 2030 3270 2045 3290
rect 2090 3270 2105 3290
rect 2030 3255 2105 3270
rect 2215 3290 2290 3305
rect 2215 3270 2230 3290
rect 2275 3270 2290 3290
rect 2215 3255 2290 3270
rect 2570 3290 2645 3305
rect 2570 3270 2585 3290
rect 2630 3270 2645 3290
rect 2570 3255 2645 3270
rect 2755 3290 2830 3305
rect 2755 3270 2770 3290
rect 2815 3270 2830 3290
rect 2755 3255 2830 3270
rect 3110 3290 3185 3305
rect 3110 3270 3125 3290
rect 3170 3270 3185 3290
rect 3110 3255 3185 3270
rect 3295 3290 3370 3305
rect 3295 3270 3310 3290
rect 3355 3270 3370 3290
rect 3295 3255 3370 3270
rect -130 2740 -55 2755
rect -130 2720 -115 2740
rect -70 2720 -55 2740
rect -130 2705 -55 2720
rect 55 2740 130 2755
rect 55 2720 70 2740
rect 115 2720 130 2740
rect 55 2705 130 2720
rect 410 2740 485 2755
rect 410 2720 425 2740
rect 470 2720 485 2740
rect 410 2705 485 2720
rect 595 2740 670 2755
rect 595 2720 610 2740
rect 655 2720 670 2740
rect 595 2705 670 2720
rect 950 2740 1025 2755
rect 950 2720 965 2740
rect 1010 2720 1025 2740
rect 950 2705 1025 2720
rect 1135 2740 1210 2755
rect 1135 2720 1150 2740
rect 1195 2720 1210 2740
rect 1135 2705 1210 2720
rect 1490 2740 1565 2755
rect 1490 2720 1505 2740
rect 1550 2720 1565 2740
rect 1490 2705 1565 2720
rect 1675 2740 1750 2755
rect 1675 2720 1690 2740
rect 1735 2720 1750 2740
rect 1675 2705 1750 2720
rect 2030 2740 2105 2755
rect 2030 2720 2045 2740
rect 2090 2720 2105 2740
rect 2030 2705 2105 2720
rect 2215 2740 2290 2755
rect 2215 2720 2230 2740
rect 2275 2720 2290 2740
rect 2215 2705 2290 2720
rect 2570 2740 2645 2755
rect 2570 2720 2585 2740
rect 2630 2720 2645 2740
rect 2570 2705 2645 2720
rect 2755 2740 2830 2755
rect 2755 2720 2770 2740
rect 2815 2720 2830 2740
rect 2755 2705 2830 2720
rect 3110 2740 3185 2755
rect 3110 2720 3125 2740
rect 3170 2720 3185 2740
rect 3110 2705 3185 2720
rect 3295 2740 3370 2755
rect 3295 2720 3310 2740
rect 3355 2720 3370 2740
rect 3295 2705 3370 2720
rect -130 2190 -55 2205
rect -130 2170 -115 2190
rect -70 2170 -55 2190
rect -130 2155 -55 2170
rect 55 2190 130 2205
rect 55 2170 70 2190
rect 115 2170 130 2190
rect 55 2155 130 2170
rect 410 2190 485 2205
rect 410 2170 425 2190
rect 470 2170 485 2190
rect 410 2155 485 2170
rect 595 2190 670 2205
rect 595 2170 610 2190
rect 655 2170 670 2190
rect 595 2155 670 2170
rect 950 2190 1025 2205
rect 950 2170 965 2190
rect 1010 2170 1025 2190
rect 950 2155 1025 2170
rect 1135 2190 1210 2205
rect 1135 2170 1150 2190
rect 1195 2170 1210 2190
rect 1135 2155 1210 2170
rect 1490 2190 1565 2205
rect 1490 2170 1505 2190
rect 1550 2170 1565 2190
rect 1490 2155 1565 2170
rect 1675 2190 1750 2205
rect 1675 2170 1690 2190
rect 1735 2170 1750 2190
rect 1675 2155 1750 2170
rect 2030 2190 2105 2205
rect 2030 2170 2045 2190
rect 2090 2170 2105 2190
rect 2030 2155 2105 2170
rect 2215 2190 2290 2205
rect 2215 2170 2230 2190
rect 2275 2170 2290 2190
rect 2215 2155 2290 2170
rect 2570 2190 2645 2205
rect 2570 2170 2585 2190
rect 2630 2170 2645 2190
rect 2570 2155 2645 2170
rect 2755 2190 2830 2205
rect 2755 2170 2770 2190
rect 2815 2170 2830 2190
rect 2755 2155 2830 2170
rect 3110 2190 3185 2205
rect 3110 2170 3125 2190
rect 3170 2170 3185 2190
rect 3110 2155 3185 2170
rect 3295 2190 3370 2205
rect 3295 2170 3310 2190
rect 3355 2170 3370 2190
rect 3295 2155 3370 2170
rect -130 1640 -55 1655
rect -130 1620 -115 1640
rect -70 1620 -55 1640
rect -130 1605 -55 1620
rect 55 1640 130 1655
rect 55 1620 70 1640
rect 115 1620 130 1640
rect 55 1605 130 1620
rect 410 1640 485 1655
rect 410 1620 425 1640
rect 470 1620 485 1640
rect 410 1605 485 1620
rect 595 1640 670 1655
rect 595 1620 610 1640
rect 655 1620 670 1640
rect 595 1605 670 1620
rect 950 1640 1025 1655
rect 950 1620 965 1640
rect 1010 1620 1025 1640
rect 950 1605 1025 1620
rect 1135 1640 1210 1655
rect 1135 1620 1150 1640
rect 1195 1620 1210 1640
rect 1135 1605 1210 1620
rect 1490 1640 1565 1655
rect 1490 1620 1505 1640
rect 1550 1620 1565 1640
rect 1490 1605 1565 1620
rect 1675 1640 1750 1655
rect 1675 1620 1690 1640
rect 1735 1620 1750 1640
rect 1675 1605 1750 1620
rect 2030 1640 2105 1655
rect 2030 1620 2045 1640
rect 2090 1620 2105 1640
rect 2030 1605 2105 1620
rect 2215 1640 2290 1655
rect 2215 1620 2230 1640
rect 2275 1620 2290 1640
rect 2215 1605 2290 1620
rect 2570 1640 2645 1655
rect 2570 1620 2585 1640
rect 2630 1620 2645 1640
rect 2570 1605 2645 1620
rect 2755 1640 2830 1655
rect 2755 1620 2770 1640
rect 2815 1620 2830 1640
rect 2755 1605 2830 1620
rect 3110 1640 3185 1655
rect 3110 1620 3125 1640
rect 3170 1620 3185 1640
rect 3110 1605 3185 1620
rect 3295 1640 3370 1655
rect 3295 1620 3310 1640
rect 3355 1620 3370 1640
rect 3295 1605 3370 1620
rect -130 1090 -55 1105
rect -130 1070 -115 1090
rect -70 1070 -55 1090
rect -130 1055 -55 1070
rect 55 1090 130 1105
rect 55 1070 70 1090
rect 115 1070 130 1090
rect 55 1055 130 1070
rect 410 1090 485 1105
rect 410 1070 425 1090
rect 470 1070 485 1090
rect 410 1055 485 1070
rect 595 1090 670 1105
rect 595 1070 610 1090
rect 655 1070 670 1090
rect 595 1055 670 1070
rect 950 1090 1025 1105
rect 950 1070 965 1090
rect 1010 1070 1025 1090
rect 950 1055 1025 1070
rect 1135 1090 1210 1105
rect 1135 1070 1150 1090
rect 1195 1070 1210 1090
rect 1135 1055 1210 1070
rect 1490 1090 1565 1105
rect 1490 1070 1505 1090
rect 1550 1070 1565 1090
rect 1490 1055 1565 1070
rect 1675 1090 1750 1105
rect 1675 1070 1690 1090
rect 1735 1070 1750 1090
rect 1675 1055 1750 1070
rect 2030 1090 2105 1105
rect 2030 1070 2045 1090
rect 2090 1070 2105 1090
rect 2030 1055 2105 1070
rect 2215 1090 2290 1105
rect 2215 1070 2230 1090
rect 2275 1070 2290 1090
rect 2215 1055 2290 1070
rect 2570 1090 2645 1105
rect 2570 1070 2585 1090
rect 2630 1070 2645 1090
rect 2570 1055 2645 1070
rect 2755 1090 2830 1105
rect 2755 1070 2770 1090
rect 2815 1070 2830 1090
rect 2755 1055 2830 1070
rect 3110 1090 3185 1105
rect 3110 1070 3125 1090
rect 3170 1070 3185 1090
rect 3110 1055 3185 1070
rect 3295 1090 3370 1105
rect 3295 1070 3310 1090
rect 3355 1070 3370 1090
rect 3295 1055 3370 1070
rect -130 540 -55 555
rect -130 520 -115 540
rect -70 520 -55 540
rect -130 505 -55 520
rect 55 540 130 555
rect 55 520 70 540
rect 115 520 130 540
rect 55 505 130 520
rect 410 540 485 555
rect 410 520 425 540
rect 470 520 485 540
rect 410 505 485 520
rect 595 540 670 555
rect 595 520 610 540
rect 655 520 670 540
rect 595 505 670 520
rect 950 540 1025 555
rect 950 520 965 540
rect 1010 520 1025 540
rect 950 505 1025 520
rect 1135 540 1210 555
rect 1135 520 1150 540
rect 1195 520 1210 540
rect 1135 505 1210 520
rect 1490 540 1565 555
rect 1490 520 1505 540
rect 1550 520 1565 540
rect 1490 505 1565 520
rect 1675 540 1750 555
rect 1675 520 1690 540
rect 1735 520 1750 540
rect 1675 505 1750 520
rect 2030 540 2105 555
rect 2030 520 2045 540
rect 2090 520 2105 540
rect 2030 505 2105 520
rect 2215 540 2290 555
rect 2215 520 2230 540
rect 2275 520 2290 540
rect 2215 505 2290 520
rect 2570 540 2645 555
rect 2570 520 2585 540
rect 2630 520 2645 540
rect 2570 505 2645 520
rect 2755 540 2830 555
rect 2755 520 2770 540
rect 2815 520 2830 540
rect 2755 505 2830 520
rect 3110 540 3185 555
rect 3110 520 3125 540
rect 3170 520 3185 540
rect 3110 505 3185 520
rect 3295 540 3370 555
rect 3295 520 3310 540
rect 3355 520 3370 540
rect 3295 505 3370 520
rect -130 410 -55 425
rect -130 390 -115 410
rect -70 390 -55 410
rect -130 375 -55 390
rect 55 410 130 425
rect 55 390 70 410
rect 115 390 130 410
rect 55 375 130 390
rect 410 410 485 425
rect 410 390 425 410
rect 470 390 485 410
rect 410 375 485 390
rect 595 410 670 425
rect 595 390 610 410
rect 655 390 670 410
rect 595 375 670 390
rect 950 410 1025 425
rect 950 390 965 410
rect 1010 390 1025 410
rect 950 375 1025 390
rect 1135 410 1210 425
rect 1135 390 1150 410
rect 1195 390 1210 410
rect 1135 375 1210 390
rect 1490 410 1565 425
rect 1490 390 1505 410
rect 1550 390 1565 410
rect 1490 375 1565 390
rect 1675 410 1750 425
rect 1675 390 1690 410
rect 1735 390 1750 410
rect 1675 375 1750 390
rect 2030 410 2105 425
rect 2030 390 2045 410
rect 2090 390 2105 410
rect 2030 375 2105 390
rect 2215 410 2290 425
rect 2215 390 2230 410
rect 2275 390 2290 410
rect 2215 375 2290 390
rect 2570 410 2645 425
rect 2570 390 2585 410
rect 2630 390 2645 410
rect 2570 375 2645 390
rect 2755 410 2830 425
rect 2755 390 2770 410
rect 2815 390 2830 410
rect 2755 375 2830 390
rect 3110 410 3185 425
rect 3110 390 3125 410
rect 3170 390 3185 410
rect 3110 375 3185 390
rect 3295 410 3370 425
rect 3295 390 3310 410
rect 3355 390 3370 410
rect 3295 375 3370 390
rect 3650 410 3725 425
rect 3650 390 3665 410
rect 3710 390 3725 410
rect 3650 375 3725 390
rect -130 -140 -55 -125
rect -130 -160 -115 -140
rect -70 -160 -55 -140
rect -130 -175 -55 -160
rect 55 -140 130 -125
rect 55 -160 70 -140
rect 115 -160 130 -140
rect 55 -175 130 -160
rect 410 -140 485 -125
rect 410 -160 425 -140
rect 470 -160 485 -140
rect 410 -175 485 -160
rect 595 -140 670 -125
rect 595 -160 610 -140
rect 655 -160 670 -140
rect 595 -175 670 -160
rect 950 -140 1025 -125
rect 950 -160 965 -140
rect 1010 -160 1025 -140
rect 950 -175 1025 -160
rect 1135 -140 1210 -125
rect 1135 -160 1150 -140
rect 1195 -160 1210 -140
rect 1135 -175 1210 -160
rect 1490 -140 1565 -125
rect 1490 -160 1505 -140
rect 1550 -160 1565 -140
rect 1490 -175 1565 -160
rect 1675 -140 1750 -125
rect 1675 -160 1690 -140
rect 1735 -160 1750 -140
rect 1675 -175 1750 -160
rect 2030 -140 2105 -125
rect 2030 -160 2045 -140
rect 2090 -160 2105 -140
rect 2030 -175 2105 -160
rect 2215 -140 2290 -125
rect 2215 -160 2230 -140
rect 2275 -160 2290 -140
rect 2215 -175 2290 -160
rect 2570 -140 2645 -125
rect 2570 -160 2585 -140
rect 2630 -160 2645 -140
rect 2570 -175 2645 -160
rect 2755 -140 2830 -125
rect 2755 -160 2770 -140
rect 2815 -160 2830 -140
rect 2755 -175 2830 -160
rect 3110 -140 3185 -125
rect 3110 -160 3125 -140
rect 3170 -160 3185 -140
rect 3110 -175 3185 -160
rect 3295 -140 3370 -125
rect 3295 -160 3310 -140
rect 3355 -160 3370 -140
rect 3295 -175 3370 -160
rect 3650 -140 3725 -125
rect 3650 -160 3665 -140
rect 3710 -160 3725 -140
rect 3650 -175 3725 -160
rect -130 -690 -55 -675
rect -130 -710 -115 -690
rect -70 -710 -55 -690
rect -130 -725 -55 -710
rect 55 -690 130 -675
rect 55 -710 70 -690
rect 115 -710 130 -690
rect 55 -725 130 -710
rect 410 -690 485 -675
rect 410 -710 425 -690
rect 470 -710 485 -690
rect 410 -725 485 -710
rect 595 -690 670 -675
rect 595 -710 610 -690
rect 655 -710 670 -690
rect 595 -725 670 -710
rect 950 -690 1025 -675
rect 950 -710 965 -690
rect 1010 -710 1025 -690
rect 950 -725 1025 -710
rect 1135 -690 1210 -675
rect 1135 -710 1150 -690
rect 1195 -710 1210 -690
rect 1135 -725 1210 -710
rect 1490 -690 1565 -675
rect 1490 -710 1505 -690
rect 1550 -710 1565 -690
rect 1490 -725 1565 -710
rect 1675 -690 1750 -675
rect 1675 -710 1690 -690
rect 1735 -710 1750 -690
rect 1675 -725 1750 -710
rect 2030 -690 2105 -675
rect 2030 -710 2045 -690
rect 2090 -710 2105 -690
rect 2030 -725 2105 -710
rect 2215 -690 2290 -675
rect 2215 -710 2230 -690
rect 2275 -710 2290 -690
rect 2215 -725 2290 -710
rect 2570 -690 2645 -675
rect 2570 -710 2585 -690
rect 2630 -710 2645 -690
rect 2570 -725 2645 -710
rect 2755 -690 2830 -675
rect 2755 -710 2770 -690
rect 2815 -710 2830 -690
rect 2755 -725 2830 -710
rect 3110 -690 3185 -675
rect 3110 -710 3125 -690
rect 3170 -710 3185 -690
rect 3110 -725 3185 -710
rect 3295 -690 3370 -675
rect 3295 -710 3310 -690
rect 3355 -710 3370 -690
rect 3295 -725 3370 -710
rect 3650 -690 3725 -675
rect 3650 -710 3665 -690
rect 3710 -710 3725 -690
rect 3650 -725 3725 -710
rect -130 -1240 -55 -1225
rect -130 -1260 -115 -1240
rect -70 -1260 -55 -1240
rect -130 -1275 -55 -1260
rect 55 -1240 130 -1225
rect 55 -1260 70 -1240
rect 115 -1260 130 -1240
rect 55 -1275 130 -1260
rect 410 -1240 485 -1225
rect 410 -1260 425 -1240
rect 470 -1260 485 -1240
rect 410 -1275 485 -1260
rect 595 -1240 670 -1225
rect 595 -1260 610 -1240
rect 655 -1260 670 -1240
rect 595 -1275 670 -1260
rect 950 -1240 1025 -1225
rect 950 -1260 965 -1240
rect 1010 -1260 1025 -1240
rect 950 -1275 1025 -1260
rect 1135 -1240 1210 -1225
rect 1135 -1260 1150 -1240
rect 1195 -1260 1210 -1240
rect 1135 -1275 1210 -1260
rect 1490 -1240 1565 -1225
rect 1490 -1260 1505 -1240
rect 1550 -1260 1565 -1240
rect 1490 -1275 1565 -1260
rect 1675 -1240 1750 -1225
rect 1675 -1260 1690 -1240
rect 1735 -1260 1750 -1240
rect 1675 -1275 1750 -1260
rect 2030 -1240 2105 -1225
rect 2030 -1260 2045 -1240
rect 2090 -1260 2105 -1240
rect 2030 -1275 2105 -1260
rect 2215 -1240 2290 -1225
rect 2215 -1260 2230 -1240
rect 2275 -1260 2290 -1240
rect 2215 -1275 2290 -1260
rect 2570 -1240 2645 -1225
rect 2570 -1260 2585 -1240
rect 2630 -1260 2645 -1240
rect 2570 -1275 2645 -1260
rect 2755 -1240 2830 -1225
rect 2755 -1260 2770 -1240
rect 2815 -1260 2830 -1240
rect 2755 -1275 2830 -1260
rect 3110 -1240 3185 -1225
rect 3110 -1260 3125 -1240
rect 3170 -1260 3185 -1240
rect 3110 -1275 3185 -1260
rect 3295 -1240 3370 -1225
rect 3295 -1260 3310 -1240
rect 3355 -1260 3370 -1240
rect 3295 -1275 3370 -1260
rect 3650 -1240 3725 -1225
rect 3650 -1260 3665 -1240
rect 3710 -1260 3725 -1240
rect 3650 -1275 3725 -1260
rect -130 -1790 -55 -1775
rect -130 -1810 -115 -1790
rect -70 -1810 -55 -1790
rect -130 -1825 -55 -1810
rect 55 -1790 130 -1775
rect 55 -1810 70 -1790
rect 115 -1810 130 -1790
rect 55 -1825 130 -1810
rect 410 -1790 485 -1775
rect 410 -1810 425 -1790
rect 470 -1810 485 -1790
rect 410 -1825 485 -1810
rect 595 -1790 670 -1775
rect 595 -1810 610 -1790
rect 655 -1810 670 -1790
rect 595 -1825 670 -1810
rect 950 -1790 1025 -1775
rect 950 -1810 965 -1790
rect 1010 -1810 1025 -1790
rect 950 -1825 1025 -1810
rect 1135 -1790 1210 -1775
rect 1135 -1810 1150 -1790
rect 1195 -1810 1210 -1790
rect 1135 -1825 1210 -1810
rect 1490 -1790 1565 -1775
rect 1490 -1810 1505 -1790
rect 1550 -1810 1565 -1790
rect 1490 -1825 1565 -1810
rect 1675 -1790 1750 -1775
rect 1675 -1810 1690 -1790
rect 1735 -1810 1750 -1790
rect 1675 -1825 1750 -1810
rect 2030 -1790 2105 -1775
rect 2030 -1810 2045 -1790
rect 2090 -1810 2105 -1790
rect 2030 -1825 2105 -1810
rect 2215 -1790 2290 -1775
rect 2215 -1810 2230 -1790
rect 2275 -1810 2290 -1790
rect 2215 -1825 2290 -1810
rect 2570 -1790 2645 -1775
rect 2570 -1810 2585 -1790
rect 2630 -1810 2645 -1790
rect 2570 -1825 2645 -1810
rect 2755 -1790 2830 -1775
rect 2755 -1810 2770 -1790
rect 2815 -1810 2830 -1790
rect 2755 -1825 2830 -1810
rect 3110 -1790 3185 -1775
rect 3110 -1810 3125 -1790
rect 3170 -1810 3185 -1790
rect 3110 -1825 3185 -1810
rect 3295 -1790 3370 -1775
rect 3295 -1810 3310 -1790
rect 3355 -1810 3370 -1790
rect 3295 -1825 3370 -1810
rect 3650 -1790 3725 -1775
rect 3650 -1810 3665 -1790
rect 3710 -1810 3725 -1790
rect 3650 -1825 3725 -1810
rect -130 -2340 -55 -2325
rect -130 -2360 -115 -2340
rect -70 -2360 -55 -2340
rect -130 -2375 -55 -2360
rect 55 -2340 130 -2325
rect 55 -2360 70 -2340
rect 115 -2360 130 -2340
rect 55 -2375 130 -2360
rect 410 -2340 485 -2325
rect 410 -2360 425 -2340
rect 470 -2360 485 -2340
rect 410 -2375 485 -2360
rect 595 -2340 670 -2325
rect 595 -2360 610 -2340
rect 655 -2360 670 -2340
rect 595 -2375 670 -2360
rect 950 -2340 1025 -2325
rect 950 -2360 965 -2340
rect 1010 -2360 1025 -2340
rect 950 -2375 1025 -2360
rect 1135 -2340 1210 -2325
rect 1135 -2360 1150 -2340
rect 1195 -2360 1210 -2340
rect 1135 -2375 1210 -2360
rect 1490 -2340 1565 -2325
rect 1490 -2360 1505 -2340
rect 1550 -2360 1565 -2340
rect 1490 -2375 1565 -2360
rect 1675 -2340 1750 -2325
rect 1675 -2360 1690 -2340
rect 1735 -2360 1750 -2340
rect 1675 -2375 1750 -2360
rect 2030 -2340 2105 -2325
rect 2030 -2360 2045 -2340
rect 2090 -2360 2105 -2340
rect 2030 -2375 2105 -2360
rect 2215 -2340 2290 -2325
rect 2215 -2360 2230 -2340
rect 2275 -2360 2290 -2340
rect 2215 -2375 2290 -2360
rect 2570 -2340 2645 -2325
rect 2570 -2360 2585 -2340
rect 2630 -2360 2645 -2340
rect 2570 -2375 2645 -2360
rect 2755 -2340 2830 -2325
rect 2755 -2360 2770 -2340
rect 2815 -2360 2830 -2340
rect 2755 -2375 2830 -2360
rect 3110 -2340 3185 -2325
rect 3110 -2360 3125 -2340
rect 3170 -2360 3185 -2340
rect 3110 -2375 3185 -2360
rect 3295 -2340 3370 -2325
rect 3295 -2360 3310 -2340
rect 3355 -2360 3370 -2340
rect 3295 -2375 3370 -2360
rect 3650 -2340 3725 -2325
rect 3650 -2360 3665 -2340
rect 3710 -2360 3725 -2340
rect 3650 -2375 3725 -2360
rect -130 -2425 -55 -2410
rect -130 -2445 -115 -2425
rect -70 -2445 -55 -2425
rect -130 -2460 -55 -2445
rect 55 -2425 130 -2410
rect 55 -2445 70 -2425
rect 115 -2445 130 -2425
rect 55 -2460 130 -2445
rect 410 -2425 485 -2410
rect 410 -2445 425 -2425
rect 470 -2445 485 -2425
rect 410 -2460 485 -2445
rect 595 -2425 670 -2410
rect 595 -2445 610 -2425
rect 655 -2445 670 -2425
rect 595 -2460 670 -2445
rect 950 -2425 1025 -2410
rect 950 -2445 965 -2425
rect 1010 -2445 1025 -2425
rect 950 -2460 1025 -2445
rect 1135 -2425 1210 -2410
rect 1135 -2445 1150 -2425
rect 1195 -2445 1210 -2425
rect 1135 -2460 1210 -2445
rect 1490 -2425 1565 -2410
rect 1490 -2445 1505 -2425
rect 1550 -2445 1565 -2425
rect 1490 -2460 1565 -2445
rect 1675 -2425 1750 -2410
rect 1675 -2445 1690 -2425
rect 1735 -2445 1750 -2425
rect 1675 -2460 1750 -2445
rect 2030 -2425 2105 -2410
rect 2030 -2445 2045 -2425
rect 2090 -2445 2105 -2425
rect 2030 -2460 2105 -2445
rect 2215 -2425 2290 -2410
rect 2215 -2445 2230 -2425
rect 2275 -2445 2290 -2425
rect 2215 -2460 2290 -2445
rect 2570 -2425 2645 -2410
rect 2570 -2445 2585 -2425
rect 2630 -2445 2645 -2425
rect 2570 -2460 2645 -2445
rect 2755 -2425 2830 -2410
rect 2755 -2445 2770 -2425
rect 2815 -2445 2830 -2425
rect 2755 -2460 2830 -2445
rect 3110 -2425 3185 -2410
rect 3110 -2445 3125 -2425
rect 3170 -2445 3185 -2425
rect 3110 -2460 3185 -2445
rect 3295 -2425 3370 -2410
rect 3295 -2445 3310 -2425
rect 3355 -2445 3370 -2425
rect 3295 -2460 3370 -2445
rect 3650 -2425 3725 -2410
rect 3650 -2445 3665 -2425
rect 3710 -2445 3725 -2425
rect 3650 -2460 3725 -2445
rect -130 -2975 -55 -2960
rect -130 -2995 -115 -2975
rect -70 -2995 -55 -2975
rect -130 -3010 -55 -2995
rect 55 -2975 130 -2960
rect 55 -2995 70 -2975
rect 115 -2995 130 -2975
rect 55 -3010 130 -2995
rect 410 -2975 485 -2960
rect 410 -2995 425 -2975
rect 470 -2995 485 -2975
rect 410 -3010 485 -2995
rect 595 -2975 670 -2960
rect 595 -2995 610 -2975
rect 655 -2995 670 -2975
rect 595 -3010 670 -2995
rect 950 -2975 1025 -2960
rect 950 -2995 965 -2975
rect 1010 -2995 1025 -2975
rect 950 -3010 1025 -2995
rect 1135 -2975 1210 -2960
rect 1135 -2995 1150 -2975
rect 1195 -2995 1210 -2975
rect 1135 -3010 1210 -2995
rect 1490 -2975 1565 -2960
rect 1490 -2995 1505 -2975
rect 1550 -2995 1565 -2975
rect 1490 -3010 1565 -2995
rect 1675 -2975 1750 -2960
rect 1675 -2995 1690 -2975
rect 1735 -2995 1750 -2975
rect 1675 -3010 1750 -2995
rect 2030 -2975 2105 -2960
rect 2030 -2995 2045 -2975
rect 2090 -2995 2105 -2975
rect 2030 -3010 2105 -2995
rect 2215 -2975 2290 -2960
rect 2215 -2995 2230 -2975
rect 2275 -2995 2290 -2975
rect 2215 -3010 2290 -2995
rect 2570 -2975 2645 -2960
rect 2570 -2995 2585 -2975
rect 2630 -2995 2645 -2975
rect 2570 -3010 2645 -2995
rect 2755 -2975 2830 -2960
rect 2755 -2995 2770 -2975
rect 2815 -2995 2830 -2975
rect 2755 -3010 2830 -2995
rect 3110 -2975 3185 -2960
rect 3110 -2995 3125 -2975
rect 3170 -2995 3185 -2975
rect 3110 -3010 3185 -2995
rect 3295 -2975 3370 -2960
rect 3295 -2995 3310 -2975
rect 3355 -2995 3370 -2975
rect 3295 -3010 3370 -2995
rect 3650 -2975 3725 -2960
rect 3650 -2995 3665 -2975
rect 3710 -2995 3725 -2975
rect 3650 -3010 3725 -2995
rect -130 -3525 -55 -3510
rect -130 -3545 -115 -3525
rect -70 -3545 -55 -3525
rect -130 -3560 -55 -3545
rect 55 -3525 130 -3510
rect 55 -3545 70 -3525
rect 115 -3545 130 -3525
rect 55 -3560 130 -3545
rect 410 -3525 485 -3510
rect 410 -3545 425 -3525
rect 470 -3545 485 -3525
rect 410 -3560 485 -3545
rect 595 -3525 670 -3510
rect 595 -3545 610 -3525
rect 655 -3545 670 -3525
rect 595 -3560 670 -3545
rect 950 -3525 1025 -3510
rect 950 -3545 965 -3525
rect 1010 -3545 1025 -3525
rect 950 -3560 1025 -3545
rect 1135 -3525 1210 -3510
rect 1135 -3545 1150 -3525
rect 1195 -3545 1210 -3525
rect 1135 -3560 1210 -3545
rect 1490 -3525 1565 -3510
rect 1490 -3545 1505 -3525
rect 1550 -3545 1565 -3525
rect 1490 -3560 1565 -3545
rect 1675 -3525 1750 -3510
rect 1675 -3545 1690 -3525
rect 1735 -3545 1750 -3525
rect 1675 -3560 1750 -3545
rect 2030 -3525 2105 -3510
rect 2030 -3545 2045 -3525
rect 2090 -3545 2105 -3525
rect 2030 -3560 2105 -3545
rect 2215 -3525 2290 -3510
rect 2215 -3545 2230 -3525
rect 2275 -3545 2290 -3525
rect 2215 -3560 2290 -3545
rect 2570 -3525 2645 -3510
rect 2570 -3545 2585 -3525
rect 2630 -3545 2645 -3525
rect 2570 -3560 2645 -3545
rect 2755 -3525 2830 -3510
rect 2755 -3545 2770 -3525
rect 2815 -3545 2830 -3525
rect 2755 -3560 2830 -3545
rect 3110 -3525 3185 -3510
rect 3110 -3545 3125 -3525
rect 3170 -3545 3185 -3525
rect 3110 -3560 3185 -3545
rect 3295 -3525 3370 -3510
rect 3295 -3545 3310 -3525
rect 3355 -3545 3370 -3525
rect 3295 -3560 3370 -3545
rect 3650 -3525 3725 -3510
rect 3650 -3545 3665 -3525
rect 3710 -3545 3725 -3525
rect 3650 -3560 3725 -3545
rect -130 -4075 -55 -4060
rect -130 -4095 -115 -4075
rect -70 -4095 -55 -4075
rect -130 -4110 -55 -4095
rect 55 -4075 130 -4060
rect 55 -4095 70 -4075
rect 115 -4095 130 -4075
rect 55 -4110 130 -4095
rect 410 -4075 485 -4060
rect 410 -4095 425 -4075
rect 470 -4095 485 -4075
rect 410 -4110 485 -4095
rect 595 -4075 670 -4060
rect 595 -4095 610 -4075
rect 655 -4095 670 -4075
rect 595 -4110 670 -4095
rect 950 -4075 1025 -4060
rect 950 -4095 965 -4075
rect 1010 -4095 1025 -4075
rect 950 -4110 1025 -4095
rect 1135 -4075 1210 -4060
rect 1135 -4095 1150 -4075
rect 1195 -4095 1210 -4075
rect 1135 -4110 1210 -4095
rect 1490 -4075 1565 -4060
rect 1490 -4095 1505 -4075
rect 1550 -4095 1565 -4075
rect 1490 -4110 1565 -4095
rect 1675 -4075 1750 -4060
rect 1675 -4095 1690 -4075
rect 1735 -4095 1750 -4075
rect 1675 -4110 1750 -4095
rect 2030 -4075 2105 -4060
rect 2030 -4095 2045 -4075
rect 2090 -4095 2105 -4075
rect 2030 -4110 2105 -4095
rect 2215 -4075 2290 -4060
rect 2215 -4095 2230 -4075
rect 2275 -4095 2290 -4075
rect 2215 -4110 2290 -4095
rect 2570 -4075 2645 -4060
rect 2570 -4095 2585 -4075
rect 2630 -4095 2645 -4075
rect 2570 -4110 2645 -4095
rect 2755 -4075 2830 -4060
rect 2755 -4095 2770 -4075
rect 2815 -4095 2830 -4075
rect 2755 -4110 2830 -4095
rect 3110 -4075 3185 -4060
rect 3110 -4095 3125 -4075
rect 3170 -4095 3185 -4075
rect 3110 -4110 3185 -4095
rect 3295 -4075 3370 -4060
rect 3295 -4095 3310 -4075
rect 3355 -4095 3370 -4075
rect 3295 -4110 3370 -4095
rect 3650 -4075 3725 -4060
rect 3650 -4095 3665 -4075
rect 3710 -4095 3725 -4075
rect 3650 -4110 3725 -4095
rect -130 -4625 -55 -4610
rect -130 -4645 -115 -4625
rect -70 -4645 -55 -4625
rect -130 -4660 -55 -4645
rect 55 -4625 130 -4610
rect 55 -4645 70 -4625
rect 115 -4645 130 -4625
rect 55 -4660 130 -4645
rect 410 -4625 485 -4610
rect 410 -4645 425 -4625
rect 470 -4645 485 -4625
rect 410 -4660 485 -4645
rect 595 -4625 670 -4610
rect 595 -4645 610 -4625
rect 655 -4645 670 -4625
rect 595 -4660 670 -4645
rect 950 -4625 1025 -4610
rect 950 -4645 965 -4625
rect 1010 -4645 1025 -4625
rect 950 -4660 1025 -4645
rect 1135 -4625 1210 -4610
rect 1135 -4645 1150 -4625
rect 1195 -4645 1210 -4625
rect 1135 -4660 1210 -4645
rect 1490 -4625 1565 -4610
rect 1490 -4645 1505 -4625
rect 1550 -4645 1565 -4625
rect 1490 -4660 1565 -4645
rect 1675 -4625 1750 -4610
rect 1675 -4645 1690 -4625
rect 1735 -4645 1750 -4625
rect 1675 -4660 1750 -4645
rect 2030 -4625 2105 -4610
rect 2030 -4645 2045 -4625
rect 2090 -4645 2105 -4625
rect 2030 -4660 2105 -4645
rect 2215 -4625 2290 -4610
rect 2215 -4645 2230 -4625
rect 2275 -4645 2290 -4625
rect 2215 -4660 2290 -4645
rect 2570 -4625 2645 -4610
rect 2570 -4645 2585 -4625
rect 2630 -4645 2645 -4625
rect 2570 -4660 2645 -4645
rect 2755 -4625 2830 -4610
rect 2755 -4645 2770 -4625
rect 2815 -4645 2830 -4625
rect 2755 -4660 2830 -4645
rect 3110 -4625 3185 -4610
rect 3110 -4645 3125 -4625
rect 3170 -4645 3185 -4625
rect 3110 -4660 3185 -4645
rect 3295 -4625 3370 -4610
rect 3295 -4645 3310 -4625
rect 3355 -4645 3370 -4625
rect 3295 -4660 3370 -4645
rect 3650 -4625 3725 -4610
rect 3650 -4645 3665 -4625
rect 3710 -4645 3725 -4625
rect 3650 -4660 3725 -4645
rect -130 -5175 -55 -5160
rect -130 -5195 -115 -5175
rect -70 -5195 -55 -5175
rect -130 -5210 -55 -5195
rect 55 -5175 130 -5160
rect 55 -5195 70 -5175
rect 115 -5195 130 -5175
rect 55 -5210 130 -5195
rect 410 -5175 485 -5160
rect 410 -5195 425 -5175
rect 470 -5195 485 -5175
rect 410 -5210 485 -5195
rect 595 -5175 670 -5160
rect 595 -5195 610 -5175
rect 655 -5195 670 -5175
rect 595 -5210 670 -5195
rect 950 -5175 1025 -5160
rect 950 -5195 965 -5175
rect 1010 -5195 1025 -5175
rect 950 -5210 1025 -5195
rect 1135 -5175 1210 -5160
rect 1135 -5195 1150 -5175
rect 1195 -5195 1210 -5175
rect 1135 -5210 1210 -5195
rect 1490 -5175 1565 -5160
rect 1490 -5195 1505 -5175
rect 1550 -5195 1565 -5175
rect 1490 -5210 1565 -5195
rect 1675 -5175 1750 -5160
rect 1675 -5195 1690 -5175
rect 1735 -5195 1750 -5175
rect 1675 -5210 1750 -5195
rect 2030 -5175 2105 -5160
rect 2030 -5195 2045 -5175
rect 2090 -5195 2105 -5175
rect 2030 -5210 2105 -5195
rect 2215 -5175 2290 -5160
rect 2215 -5195 2230 -5175
rect 2275 -5195 2290 -5175
rect 2215 -5210 2290 -5195
rect 2570 -5175 2645 -5160
rect 2570 -5195 2585 -5175
rect 2630 -5195 2645 -5175
rect 2570 -5210 2645 -5195
rect 2755 -5175 2830 -5160
rect 2755 -5195 2770 -5175
rect 2815 -5195 2830 -5175
rect 2755 -5210 2830 -5195
rect 3110 -5175 3185 -5160
rect 3110 -5195 3125 -5175
rect 3170 -5195 3185 -5175
rect 3110 -5210 3185 -5195
rect 3295 -5175 3370 -5160
rect 3295 -5195 3310 -5175
rect 3355 -5195 3370 -5175
rect 3295 -5210 3370 -5195
rect 3650 -5175 3725 -5160
rect 3650 -5195 3665 -5175
rect 3710 -5195 3725 -5175
rect 3650 -5210 3725 -5195
rect -130 -5330 -55 -5315
rect -130 -5350 -115 -5330
rect -70 -5350 -55 -5330
rect -130 -5365 -55 -5350
rect 55 -5330 130 -5315
rect 55 -5350 70 -5330
rect 115 -5350 130 -5330
rect 55 -5365 130 -5350
rect 410 -5330 485 -5315
rect 410 -5350 425 -5330
rect 470 -5350 485 -5330
rect 410 -5365 485 -5350
rect 595 -5330 670 -5315
rect 595 -5350 610 -5330
rect 655 -5350 670 -5330
rect 595 -5365 670 -5350
rect 950 -5330 1025 -5315
rect 950 -5350 965 -5330
rect 1010 -5350 1025 -5330
rect 950 -5365 1025 -5350
rect 1135 -5330 1210 -5315
rect 1135 -5350 1150 -5330
rect 1195 -5350 1210 -5330
rect 1135 -5365 1210 -5350
rect 1490 -5330 1565 -5315
rect 1490 -5350 1505 -5330
rect 1550 -5350 1565 -5330
rect 1490 -5365 1565 -5350
rect 1675 -5330 1750 -5315
rect 1675 -5350 1690 -5330
rect 1735 -5350 1750 -5330
rect 1675 -5365 1750 -5350
rect 2030 -5330 2105 -5315
rect 2030 -5350 2045 -5330
rect 2090 -5350 2105 -5330
rect 2030 -5365 2105 -5350
rect 2215 -5330 2290 -5315
rect 2215 -5350 2230 -5330
rect 2275 -5350 2290 -5330
rect 2215 -5365 2290 -5350
rect 2570 -5330 2645 -5315
rect 2570 -5350 2585 -5330
rect 2630 -5350 2645 -5330
rect 2570 -5365 2645 -5350
rect 2755 -5330 2830 -5315
rect 2755 -5350 2770 -5330
rect 2815 -5350 2830 -5330
rect 2755 -5365 2830 -5350
rect 3110 -5330 3185 -5315
rect 3110 -5350 3125 -5330
rect 3170 -5350 3185 -5330
rect 3110 -5365 3185 -5350
rect 3295 -5330 3370 -5315
rect 3295 -5350 3310 -5330
rect 3355 -5350 3370 -5330
rect 3295 -5365 3370 -5350
rect -130 -5880 -55 -5865
rect -130 -5900 -115 -5880
rect -70 -5900 -55 -5880
rect -130 -5915 -55 -5900
rect 55 -5880 130 -5865
rect 55 -5900 70 -5880
rect 115 -5900 130 -5880
rect 55 -5915 130 -5900
rect 410 -5880 485 -5865
rect 410 -5900 425 -5880
rect 470 -5900 485 -5880
rect 410 -5915 485 -5900
rect 595 -5880 670 -5865
rect 595 -5900 610 -5880
rect 655 -5900 670 -5880
rect 595 -5915 670 -5900
rect 950 -5880 1025 -5865
rect 950 -5900 965 -5880
rect 1010 -5900 1025 -5880
rect 950 -5915 1025 -5900
rect 1135 -5880 1210 -5865
rect 1135 -5900 1150 -5880
rect 1195 -5900 1210 -5880
rect 1135 -5915 1210 -5900
rect 1490 -5880 1565 -5865
rect 1490 -5900 1505 -5880
rect 1550 -5900 1565 -5880
rect 1490 -5915 1565 -5900
rect 1675 -5880 1750 -5865
rect 1675 -5900 1690 -5880
rect 1735 -5900 1750 -5880
rect 1675 -5915 1750 -5900
rect 2030 -5880 2105 -5865
rect 2030 -5900 2045 -5880
rect 2090 -5900 2105 -5880
rect 2030 -5915 2105 -5900
rect 2215 -5880 2290 -5865
rect 2215 -5900 2230 -5880
rect 2275 -5900 2290 -5880
rect 2215 -5915 2290 -5900
rect 2570 -5880 2645 -5865
rect 2570 -5900 2585 -5880
rect 2630 -5900 2645 -5880
rect 2570 -5915 2645 -5900
rect 2755 -5880 2830 -5865
rect 2755 -5900 2770 -5880
rect 2815 -5900 2830 -5880
rect 2755 -5915 2830 -5900
rect 3110 -5880 3185 -5865
rect 3110 -5900 3125 -5880
rect 3170 -5900 3185 -5880
rect 3110 -5915 3185 -5900
rect 3295 -5880 3370 -5865
rect 3295 -5900 3310 -5880
rect 3355 -5900 3370 -5880
rect 3295 -5915 3370 -5900
rect -130 -6430 -55 -6415
rect -130 -6450 -115 -6430
rect -70 -6450 -55 -6430
rect -130 -6465 -55 -6450
rect 55 -6430 130 -6415
rect 55 -6450 70 -6430
rect 115 -6450 130 -6430
rect 55 -6465 130 -6450
rect 410 -6430 485 -6415
rect 410 -6450 425 -6430
rect 470 -6450 485 -6430
rect 410 -6465 485 -6450
rect 595 -6430 670 -6415
rect 595 -6450 610 -6430
rect 655 -6450 670 -6430
rect 595 -6465 670 -6450
rect 950 -6430 1025 -6415
rect 950 -6450 965 -6430
rect 1010 -6450 1025 -6430
rect 950 -6465 1025 -6450
rect 1135 -6430 1210 -6415
rect 1135 -6450 1150 -6430
rect 1195 -6450 1210 -6430
rect 1135 -6465 1210 -6450
rect 1490 -6430 1565 -6415
rect 1490 -6450 1505 -6430
rect 1550 -6450 1565 -6430
rect 1490 -6465 1565 -6450
rect 1675 -6430 1750 -6415
rect 1675 -6450 1690 -6430
rect 1735 -6450 1750 -6430
rect 1675 -6465 1750 -6450
rect 2030 -6430 2105 -6415
rect 2030 -6450 2045 -6430
rect 2090 -6450 2105 -6430
rect 2030 -6465 2105 -6450
rect 2215 -6430 2290 -6415
rect 2215 -6450 2230 -6430
rect 2275 -6450 2290 -6430
rect 2215 -6465 2290 -6450
rect 2570 -6430 2645 -6415
rect 2570 -6450 2585 -6430
rect 2630 -6450 2645 -6430
rect 2570 -6465 2645 -6450
rect 2755 -6430 2830 -6415
rect 2755 -6450 2770 -6430
rect 2815 -6450 2830 -6430
rect 2755 -6465 2830 -6450
rect 3110 -6430 3185 -6415
rect 3110 -6450 3125 -6430
rect 3170 -6450 3185 -6430
rect 3110 -6465 3185 -6450
rect 3295 -6430 3370 -6415
rect 3295 -6450 3310 -6430
rect 3355 -6450 3370 -6430
rect 3295 -6465 3370 -6450
rect -130 -6980 -55 -6965
rect -130 -7000 -115 -6980
rect -70 -7000 -55 -6980
rect -130 -7015 -55 -7000
rect 55 -6980 130 -6965
rect 55 -7000 70 -6980
rect 115 -7000 130 -6980
rect 55 -7015 130 -7000
rect 410 -6980 485 -6965
rect 410 -7000 425 -6980
rect 470 -7000 485 -6980
rect 410 -7015 485 -7000
rect 595 -6980 670 -6965
rect 595 -7000 610 -6980
rect 655 -7000 670 -6980
rect 595 -7015 670 -7000
rect 950 -6980 1025 -6965
rect 950 -7000 965 -6980
rect 1010 -7000 1025 -6980
rect 950 -7015 1025 -7000
rect 1135 -6980 1210 -6965
rect 1135 -7000 1150 -6980
rect 1195 -7000 1210 -6980
rect 1135 -7015 1210 -7000
rect 1490 -6980 1565 -6965
rect 1490 -7000 1505 -6980
rect 1550 -7000 1565 -6980
rect 1490 -7015 1565 -7000
rect 1675 -6980 1750 -6965
rect 1675 -7000 1690 -6980
rect 1735 -7000 1750 -6980
rect 1675 -7015 1750 -7000
rect 2030 -6980 2105 -6965
rect 2030 -7000 2045 -6980
rect 2090 -7000 2105 -6980
rect 2030 -7015 2105 -7000
rect 2215 -6980 2290 -6965
rect 2215 -7000 2230 -6980
rect 2275 -7000 2290 -6980
rect 2215 -7015 2290 -7000
rect 2570 -6980 2645 -6965
rect 2570 -7000 2585 -6980
rect 2630 -7000 2645 -6980
rect 2570 -7015 2645 -7000
rect 2755 -6980 2830 -6965
rect 2755 -7000 2770 -6980
rect 2815 -7000 2830 -6980
rect 2755 -7015 2830 -7000
rect 3110 -6980 3185 -6965
rect 3110 -7000 3125 -6980
rect 3170 -7000 3185 -6980
rect 3110 -7015 3185 -7000
rect 3295 -6980 3370 -6965
rect 3295 -7000 3310 -6980
rect 3355 -7000 3370 -6980
rect 3295 -7015 3370 -7000
rect -130 -7530 -55 -7515
rect -130 -7550 -115 -7530
rect -70 -7550 -55 -7530
rect -130 -7565 -55 -7550
rect 55 -7530 130 -7515
rect 55 -7550 70 -7530
rect 115 -7550 130 -7530
rect 55 -7565 130 -7550
rect 410 -7530 485 -7515
rect 410 -7550 425 -7530
rect 470 -7550 485 -7530
rect 410 -7565 485 -7550
rect 595 -7530 670 -7515
rect 595 -7550 610 -7530
rect 655 -7550 670 -7530
rect 595 -7565 670 -7550
rect 950 -7530 1025 -7515
rect 950 -7550 965 -7530
rect 1010 -7550 1025 -7530
rect 950 -7565 1025 -7550
rect 1135 -7530 1210 -7515
rect 1135 -7550 1150 -7530
rect 1195 -7550 1210 -7530
rect 1135 -7565 1210 -7550
rect 1490 -7530 1565 -7515
rect 1490 -7550 1505 -7530
rect 1550 -7550 1565 -7530
rect 1490 -7565 1565 -7550
rect 1675 -7530 1750 -7515
rect 1675 -7550 1690 -7530
rect 1735 -7550 1750 -7530
rect 1675 -7565 1750 -7550
rect 2030 -7530 2105 -7515
rect 2030 -7550 2045 -7530
rect 2090 -7550 2105 -7530
rect 2030 -7565 2105 -7550
rect 2215 -7530 2290 -7515
rect 2215 -7550 2230 -7530
rect 2275 -7550 2290 -7530
rect 2215 -7565 2290 -7550
rect 2570 -7530 2645 -7515
rect 2570 -7550 2585 -7530
rect 2630 -7550 2645 -7530
rect 2570 -7565 2645 -7550
rect 2755 -7530 2830 -7515
rect 2755 -7550 2770 -7530
rect 2815 -7550 2830 -7530
rect 2755 -7565 2830 -7550
rect 3110 -7530 3185 -7515
rect 3110 -7550 3125 -7530
rect 3170 -7550 3185 -7530
rect 3110 -7565 3185 -7550
rect 3295 -7530 3370 -7515
rect 3295 -7550 3310 -7530
rect 3355 -7550 3370 -7530
rect 3295 -7565 3370 -7550
rect -130 -8080 -55 -8065
rect -130 -8100 -115 -8080
rect -70 -8100 -55 -8080
rect -130 -8115 -55 -8100
rect 55 -8080 130 -8065
rect 55 -8100 70 -8080
rect 115 -8100 130 -8080
rect 55 -8115 130 -8100
rect 410 -8080 485 -8065
rect 410 -8100 425 -8080
rect 470 -8100 485 -8080
rect 410 -8115 485 -8100
rect 595 -8080 670 -8065
rect 595 -8100 610 -8080
rect 655 -8100 670 -8080
rect 595 -8115 670 -8100
rect 950 -8080 1025 -8065
rect 950 -8100 965 -8080
rect 1010 -8100 1025 -8080
rect 950 -8115 1025 -8100
rect 1135 -8080 1210 -8065
rect 1135 -8100 1150 -8080
rect 1195 -8100 1210 -8080
rect 1135 -8115 1210 -8100
rect 1490 -8080 1565 -8065
rect 1490 -8100 1505 -8080
rect 1550 -8100 1565 -8080
rect 1490 -8115 1565 -8100
rect 1675 -8080 1750 -8065
rect 1675 -8100 1690 -8080
rect 1735 -8100 1750 -8080
rect 1675 -8115 1750 -8100
rect 2030 -8080 2105 -8065
rect 2030 -8100 2045 -8080
rect 2090 -8100 2105 -8080
rect 2030 -8115 2105 -8100
rect 2215 -8080 2290 -8065
rect 2215 -8100 2230 -8080
rect 2275 -8100 2290 -8080
rect 2215 -8115 2290 -8100
rect 2570 -8080 2645 -8065
rect 2570 -8100 2585 -8080
rect 2630 -8100 2645 -8080
rect 2570 -8115 2645 -8100
rect 2755 -8080 2830 -8065
rect 2755 -8100 2770 -8080
rect 2815 -8100 2830 -8080
rect 2755 -8115 2830 -8100
rect 3110 -8080 3185 -8065
rect 3110 -8100 3125 -8080
rect 3170 -8100 3185 -8080
rect 3110 -8115 3185 -8100
rect 3295 -8080 3370 -8065
rect 3295 -8100 3310 -8080
rect 3355 -8100 3370 -8080
rect 3295 -8115 3370 -8100
<< ndiffc >>
rect -115 3270 -70 3290
rect 70 3270 115 3290
rect 425 3270 470 3290
rect 610 3270 655 3290
rect 965 3270 1010 3290
rect 1150 3270 1195 3290
rect 1505 3270 1550 3290
rect 1690 3270 1735 3290
rect 2045 3270 2090 3290
rect 2230 3270 2275 3290
rect 2585 3270 2630 3290
rect 2770 3270 2815 3290
rect 3125 3270 3170 3290
rect 3310 3270 3355 3290
rect -115 2720 -70 2740
rect 70 2720 115 2740
rect 425 2720 470 2740
rect 610 2720 655 2740
rect 965 2720 1010 2740
rect 1150 2720 1195 2740
rect 1505 2720 1550 2740
rect 1690 2720 1735 2740
rect 2045 2720 2090 2740
rect 2230 2720 2275 2740
rect 2585 2720 2630 2740
rect 2770 2720 2815 2740
rect 3125 2720 3170 2740
rect 3310 2720 3355 2740
rect -115 2170 -70 2190
rect 70 2170 115 2190
rect 425 2170 470 2190
rect 610 2170 655 2190
rect 965 2170 1010 2190
rect 1150 2170 1195 2190
rect 1505 2170 1550 2190
rect 1690 2170 1735 2190
rect 2045 2170 2090 2190
rect 2230 2170 2275 2190
rect 2585 2170 2630 2190
rect 2770 2170 2815 2190
rect 3125 2170 3170 2190
rect 3310 2170 3355 2190
rect -115 1620 -70 1640
rect 70 1620 115 1640
rect 425 1620 470 1640
rect 610 1620 655 1640
rect 965 1620 1010 1640
rect 1150 1620 1195 1640
rect 1505 1620 1550 1640
rect 1690 1620 1735 1640
rect 2045 1620 2090 1640
rect 2230 1620 2275 1640
rect 2585 1620 2630 1640
rect 2770 1620 2815 1640
rect 3125 1620 3170 1640
rect 3310 1620 3355 1640
rect -115 1070 -70 1090
rect 70 1070 115 1090
rect 425 1070 470 1090
rect 610 1070 655 1090
rect 965 1070 1010 1090
rect 1150 1070 1195 1090
rect 1505 1070 1550 1090
rect 1690 1070 1735 1090
rect 2045 1070 2090 1090
rect 2230 1070 2275 1090
rect 2585 1070 2630 1090
rect 2770 1070 2815 1090
rect 3125 1070 3170 1090
rect 3310 1070 3355 1090
rect -115 520 -70 540
rect 70 520 115 540
rect 425 520 470 540
rect 610 520 655 540
rect 965 520 1010 540
rect 1150 520 1195 540
rect 1505 520 1550 540
rect 1690 520 1735 540
rect 2045 520 2090 540
rect 2230 520 2275 540
rect 2585 520 2630 540
rect 2770 520 2815 540
rect 3125 520 3170 540
rect 3310 520 3355 540
rect -115 390 -70 410
rect 70 390 115 410
rect 425 390 470 410
rect 610 390 655 410
rect 965 390 1010 410
rect 1150 390 1195 410
rect 1505 390 1550 410
rect 1690 390 1735 410
rect 2045 390 2090 410
rect 2230 390 2275 410
rect 2585 390 2630 410
rect 2770 390 2815 410
rect 3125 390 3170 410
rect 3310 390 3355 410
rect 3665 390 3710 410
rect -115 -160 -70 -140
rect 70 -160 115 -140
rect 425 -160 470 -140
rect 610 -160 655 -140
rect 965 -160 1010 -140
rect 1150 -160 1195 -140
rect 1505 -160 1550 -140
rect 1690 -160 1735 -140
rect 2045 -160 2090 -140
rect 2230 -160 2275 -140
rect 2585 -160 2630 -140
rect 2770 -160 2815 -140
rect 3125 -160 3170 -140
rect 3310 -160 3355 -140
rect 3665 -160 3710 -140
rect -115 -710 -70 -690
rect 70 -710 115 -690
rect 425 -710 470 -690
rect 610 -710 655 -690
rect 965 -710 1010 -690
rect 1150 -710 1195 -690
rect 1505 -710 1550 -690
rect 1690 -710 1735 -690
rect 2045 -710 2090 -690
rect 2230 -710 2275 -690
rect 2585 -710 2630 -690
rect 2770 -710 2815 -690
rect 3125 -710 3170 -690
rect 3310 -710 3355 -690
rect 3665 -710 3710 -690
rect -115 -1260 -70 -1240
rect 70 -1260 115 -1240
rect 425 -1260 470 -1240
rect 610 -1260 655 -1240
rect 965 -1260 1010 -1240
rect 1150 -1260 1195 -1240
rect 1505 -1260 1550 -1240
rect 1690 -1260 1735 -1240
rect 2045 -1260 2090 -1240
rect 2230 -1260 2275 -1240
rect 2585 -1260 2630 -1240
rect 2770 -1260 2815 -1240
rect 3125 -1260 3170 -1240
rect 3310 -1260 3355 -1240
rect 3665 -1260 3710 -1240
rect -115 -1810 -70 -1790
rect 70 -1810 115 -1790
rect 425 -1810 470 -1790
rect 610 -1810 655 -1790
rect 965 -1810 1010 -1790
rect 1150 -1810 1195 -1790
rect 1505 -1810 1550 -1790
rect 1690 -1810 1735 -1790
rect 2045 -1810 2090 -1790
rect 2230 -1810 2275 -1790
rect 2585 -1810 2630 -1790
rect 2770 -1810 2815 -1790
rect 3125 -1810 3170 -1790
rect 3310 -1810 3355 -1790
rect 3665 -1810 3710 -1790
rect -115 -2360 -70 -2340
rect 70 -2360 115 -2340
rect 425 -2360 470 -2340
rect 610 -2360 655 -2340
rect 965 -2360 1010 -2340
rect 1150 -2360 1195 -2340
rect 1505 -2360 1550 -2340
rect 1690 -2360 1735 -2340
rect 2045 -2360 2090 -2340
rect 2230 -2360 2275 -2340
rect 2585 -2360 2630 -2340
rect 2770 -2360 2815 -2340
rect 3125 -2360 3170 -2340
rect 3310 -2360 3355 -2340
rect 3665 -2360 3710 -2340
rect -115 -2445 -70 -2425
rect 70 -2445 115 -2425
rect 425 -2445 470 -2425
rect 610 -2445 655 -2425
rect 965 -2445 1010 -2425
rect 1150 -2445 1195 -2425
rect 1505 -2445 1550 -2425
rect 1690 -2445 1735 -2425
rect 2045 -2445 2090 -2425
rect 2230 -2445 2275 -2425
rect 2585 -2445 2630 -2425
rect 2770 -2445 2815 -2425
rect 3125 -2445 3170 -2425
rect 3310 -2445 3355 -2425
rect 3665 -2445 3710 -2425
rect -115 -2995 -70 -2975
rect 70 -2995 115 -2975
rect 425 -2995 470 -2975
rect 610 -2995 655 -2975
rect 965 -2995 1010 -2975
rect 1150 -2995 1195 -2975
rect 1505 -2995 1550 -2975
rect 1690 -2995 1735 -2975
rect 2045 -2995 2090 -2975
rect 2230 -2995 2275 -2975
rect 2585 -2995 2630 -2975
rect 2770 -2995 2815 -2975
rect 3125 -2995 3170 -2975
rect 3310 -2995 3355 -2975
rect 3665 -2995 3710 -2975
rect -115 -3545 -70 -3525
rect 70 -3545 115 -3525
rect 425 -3545 470 -3525
rect 610 -3545 655 -3525
rect 965 -3545 1010 -3525
rect 1150 -3545 1195 -3525
rect 1505 -3545 1550 -3525
rect 1690 -3545 1735 -3525
rect 2045 -3545 2090 -3525
rect 2230 -3545 2275 -3525
rect 2585 -3545 2630 -3525
rect 2770 -3545 2815 -3525
rect 3125 -3545 3170 -3525
rect 3310 -3545 3355 -3525
rect 3665 -3545 3710 -3525
rect -115 -4095 -70 -4075
rect 70 -4095 115 -4075
rect 425 -4095 470 -4075
rect 610 -4095 655 -4075
rect 965 -4095 1010 -4075
rect 1150 -4095 1195 -4075
rect 1505 -4095 1550 -4075
rect 1690 -4095 1735 -4075
rect 2045 -4095 2090 -4075
rect 2230 -4095 2275 -4075
rect 2585 -4095 2630 -4075
rect 2770 -4095 2815 -4075
rect 3125 -4095 3170 -4075
rect 3310 -4095 3355 -4075
rect 3665 -4095 3710 -4075
rect -115 -4645 -70 -4625
rect 70 -4645 115 -4625
rect 425 -4645 470 -4625
rect 610 -4645 655 -4625
rect 965 -4645 1010 -4625
rect 1150 -4645 1195 -4625
rect 1505 -4645 1550 -4625
rect 1690 -4645 1735 -4625
rect 2045 -4645 2090 -4625
rect 2230 -4645 2275 -4625
rect 2585 -4645 2630 -4625
rect 2770 -4645 2815 -4625
rect 3125 -4645 3170 -4625
rect 3310 -4645 3355 -4625
rect 3665 -4645 3710 -4625
rect -115 -5195 -70 -5175
rect 70 -5195 115 -5175
rect 425 -5195 470 -5175
rect 610 -5195 655 -5175
rect 965 -5195 1010 -5175
rect 1150 -5195 1195 -5175
rect 1505 -5195 1550 -5175
rect 1690 -5195 1735 -5175
rect 2045 -5195 2090 -5175
rect 2230 -5195 2275 -5175
rect 2585 -5195 2630 -5175
rect 2770 -5195 2815 -5175
rect 3125 -5195 3170 -5175
rect 3310 -5195 3355 -5175
rect 3665 -5195 3710 -5175
rect -115 -5350 -70 -5330
rect 70 -5350 115 -5330
rect 425 -5350 470 -5330
rect 610 -5350 655 -5330
rect 965 -5350 1010 -5330
rect 1150 -5350 1195 -5330
rect 1505 -5350 1550 -5330
rect 1690 -5350 1735 -5330
rect 2045 -5350 2090 -5330
rect 2230 -5350 2275 -5330
rect 2585 -5350 2630 -5330
rect 2770 -5350 2815 -5330
rect 3125 -5350 3170 -5330
rect 3310 -5350 3355 -5330
rect -115 -5900 -70 -5880
rect 70 -5900 115 -5880
rect 425 -5900 470 -5880
rect 610 -5900 655 -5880
rect 965 -5900 1010 -5880
rect 1150 -5900 1195 -5880
rect 1505 -5900 1550 -5880
rect 1690 -5900 1735 -5880
rect 2045 -5900 2090 -5880
rect 2230 -5900 2275 -5880
rect 2585 -5900 2630 -5880
rect 2770 -5900 2815 -5880
rect 3125 -5900 3170 -5880
rect 3310 -5900 3355 -5880
rect -115 -6450 -70 -6430
rect 70 -6450 115 -6430
rect 425 -6450 470 -6430
rect 610 -6450 655 -6430
rect 965 -6450 1010 -6430
rect 1150 -6450 1195 -6430
rect 1505 -6450 1550 -6430
rect 1690 -6450 1735 -6430
rect 2045 -6450 2090 -6430
rect 2230 -6450 2275 -6430
rect 2585 -6450 2630 -6430
rect 2770 -6450 2815 -6430
rect 3125 -6450 3170 -6430
rect 3310 -6450 3355 -6430
rect -115 -7000 -70 -6980
rect 70 -7000 115 -6980
rect 425 -7000 470 -6980
rect 610 -7000 655 -6980
rect 965 -7000 1010 -6980
rect 1150 -7000 1195 -6980
rect 1505 -7000 1550 -6980
rect 1690 -7000 1735 -6980
rect 2045 -7000 2090 -6980
rect 2230 -7000 2275 -6980
rect 2585 -7000 2630 -6980
rect 2770 -7000 2815 -6980
rect 3125 -7000 3170 -6980
rect 3310 -7000 3355 -6980
rect -115 -7550 -70 -7530
rect 70 -7550 115 -7530
rect 425 -7550 470 -7530
rect 610 -7550 655 -7530
rect 965 -7550 1010 -7530
rect 1150 -7550 1195 -7530
rect 1505 -7550 1550 -7530
rect 1690 -7550 1735 -7530
rect 2045 -7550 2090 -7530
rect 2230 -7550 2275 -7530
rect 2585 -7550 2630 -7530
rect 2770 -7550 2815 -7530
rect 3125 -7550 3170 -7530
rect 3310 -7550 3355 -7530
rect -115 -8100 -70 -8080
rect 70 -8100 115 -8080
rect 425 -8100 470 -8080
rect 610 -8100 655 -8080
rect 965 -8100 1010 -8080
rect 1150 -8100 1195 -8080
rect 1505 -8100 1550 -8080
rect 1690 -8100 1735 -8080
rect 2045 -8100 2090 -8080
rect 2230 -8100 2275 -8080
rect 2585 -8100 2630 -8080
rect 2770 -8100 2815 -8080
rect 3125 -8100 3170 -8080
rect 3310 -8100 3355 -8080
<< psubdiff >>
rect -25 1860 25 1875
rect -25 1790 -10 1860
rect 10 1790 25 1860
rect -25 1775 25 1790
rect 515 1860 565 1875
rect 515 1790 530 1860
rect 550 1790 565 1860
rect 515 1775 565 1790
rect 1055 1860 1105 1875
rect 1055 1790 1070 1860
rect 1090 1790 1105 1860
rect 1055 1775 1105 1790
rect 1595 1860 1645 1875
rect 1595 1790 1610 1860
rect 1630 1790 1645 1860
rect 1595 1775 1645 1790
rect 2135 1860 2185 1875
rect 2135 1790 2150 1860
rect 2170 1790 2185 1860
rect 2135 1775 2185 1790
rect 2675 1860 2725 1875
rect 2675 1790 2690 1860
rect 2710 1790 2725 1860
rect 2675 1775 2725 1790
rect 3215 1860 3265 1875
rect 3215 1790 3230 1860
rect 3250 1790 3265 1860
rect 3215 1775 3265 1790
rect -25 -1020 25 -1005
rect -25 -1090 -10 -1020
rect 10 -1090 25 -1020
rect -25 -1105 25 -1090
rect 515 -1020 565 -1005
rect 515 -1090 530 -1020
rect 550 -1090 565 -1020
rect 515 -1105 565 -1090
rect 1055 -1020 1105 -1005
rect 1055 -1090 1070 -1020
rect 1090 -1090 1105 -1020
rect 1055 -1105 1105 -1090
rect 1595 -1020 1645 -1005
rect 1595 -1090 1610 -1020
rect 1630 -1090 1645 -1020
rect 1595 -1105 1645 -1090
rect 2135 -1020 2185 -1005
rect 2135 -1090 2150 -1020
rect 2170 -1090 2185 -1020
rect 2135 -1105 2185 -1090
rect 2675 -1020 2725 -1005
rect 2675 -1090 2690 -1020
rect 2710 -1090 2725 -1020
rect 2675 -1105 2725 -1090
rect 3215 -1020 3265 -1005
rect 3215 -1090 3230 -1020
rect 3250 -1090 3265 -1020
rect 3215 -1105 3265 -1090
rect -25 -3855 25 -3840
rect -25 -3925 -10 -3855
rect 10 -3925 25 -3855
rect -25 -3940 25 -3925
rect 515 -3855 565 -3840
rect 515 -3925 530 -3855
rect 550 -3925 565 -3855
rect 515 -3940 565 -3925
rect 1055 -3855 1105 -3840
rect 1055 -3925 1070 -3855
rect 1090 -3925 1105 -3855
rect 1055 -3940 1105 -3925
rect 1595 -3855 1645 -3840
rect 1595 -3925 1610 -3855
rect 1630 -3925 1645 -3855
rect 1595 -3940 1645 -3925
rect 2135 -3855 2185 -3840
rect 2135 -3925 2150 -3855
rect 2170 -3925 2185 -3855
rect 2135 -3940 2185 -3925
rect 2675 -3855 2725 -3840
rect 2675 -3925 2690 -3855
rect 2710 -3925 2725 -3855
rect 2675 -3940 2725 -3925
rect 3215 -3855 3265 -3840
rect 3215 -3925 3230 -3855
rect 3250 -3925 3265 -3855
rect 3215 -3940 3265 -3925
rect -25 -6760 25 -6745
rect -25 -6830 -10 -6760
rect 10 -6830 25 -6760
rect -25 -6845 25 -6830
rect 515 -6760 565 -6745
rect 515 -6830 530 -6760
rect 550 -6830 565 -6760
rect 515 -6845 565 -6830
rect 1055 -6760 1105 -6745
rect 1055 -6830 1070 -6760
rect 1090 -6830 1105 -6760
rect 1055 -6845 1105 -6830
rect 1595 -6760 1645 -6745
rect 1595 -6830 1610 -6760
rect 1630 -6830 1645 -6760
rect 1595 -6845 1645 -6830
rect 2135 -6760 2185 -6745
rect 2135 -6830 2150 -6760
rect 2170 -6830 2185 -6760
rect 2135 -6845 2185 -6830
rect 2675 -6760 2725 -6745
rect 2675 -6830 2690 -6760
rect 2710 -6830 2725 -6760
rect 2675 -6845 2725 -6830
rect 3215 -6760 3265 -6745
rect 3215 -6830 3230 -6760
rect 3250 -6830 3265 -6760
rect 3215 -6845 3265 -6830
<< psubdiffcont >>
rect -10 1790 10 1860
rect 530 1790 550 1860
rect 1070 1790 1090 1860
rect 1610 1790 1630 1860
rect 2150 1790 2170 1860
rect 2690 1790 2710 1860
rect 3230 1790 3250 1860
rect -10 -1090 10 -1020
rect 530 -1090 550 -1020
rect 1070 -1090 1090 -1020
rect 1610 -1090 1630 -1020
rect 2150 -1090 2170 -1020
rect 2690 -1090 2710 -1020
rect 3230 -1090 3250 -1020
rect -10 -3925 10 -3855
rect 530 -3925 550 -3855
rect 1070 -3925 1090 -3855
rect 1610 -3925 1630 -3855
rect 2150 -3925 2170 -3855
rect 2690 -3925 2710 -3855
rect 3230 -3925 3250 -3855
rect -10 -6830 10 -6760
rect 530 -6830 550 -6760
rect 1070 -6830 1090 -6760
rect 1610 -6830 1630 -6760
rect 2150 -6830 2170 -6760
rect 2690 -6830 2710 -6760
rect 3230 -6830 3250 -6760
<< poly >>
rect -145 2755 -130 3255
rect -55 3050 -40 3255
rect -55 3040 0 3050
rect -55 3020 -30 3040
rect -10 3020 0 3040
rect -55 3010 0 3020
rect -55 2755 -40 3010
rect 40 2755 55 3255
rect 130 3050 145 3255
rect 395 3050 410 3255
rect 130 3040 185 3050
rect 130 3020 155 3040
rect 175 3020 185 3040
rect 130 3010 185 3020
rect 355 3040 410 3050
rect 355 3020 365 3040
rect 385 3020 410 3040
rect 355 3010 410 3020
rect 130 2755 145 3010
rect 395 2755 410 3010
rect 485 2755 500 3255
rect 580 2755 595 3255
rect 670 3050 685 3255
rect 935 3050 950 3255
rect 670 3040 725 3050
rect 670 3020 695 3040
rect 715 3020 725 3040
rect 670 3010 725 3020
rect 895 3040 950 3050
rect 895 3020 905 3040
rect 925 3020 950 3040
rect 895 3010 950 3020
rect 670 2755 685 3010
rect 935 2755 950 3010
rect 1025 2755 1040 3255
rect 1120 2755 1135 3255
rect 1210 3050 1225 3255
rect 1475 3050 1490 3255
rect 1210 3040 1265 3050
rect 1210 3020 1235 3040
rect 1255 3020 1265 3040
rect 1210 3010 1265 3020
rect 1435 3040 1490 3050
rect 1435 3020 1445 3040
rect 1465 3020 1490 3040
rect 1435 3010 1490 3020
rect 1210 2755 1225 3010
rect 1475 2755 1490 3010
rect 1565 2755 1580 3255
rect 1660 2755 1675 3255
rect 1750 3050 1765 3255
rect 2015 3050 2030 3255
rect 1750 3040 1805 3050
rect 1750 3020 1775 3040
rect 1795 3020 1805 3040
rect 1750 3010 1805 3020
rect 1975 3040 2030 3050
rect 1975 3020 1985 3040
rect 2005 3020 2030 3040
rect 1975 3010 2030 3020
rect 1750 2755 1765 3010
rect 2015 2755 2030 3010
rect 2105 2755 2120 3255
rect 2200 2755 2215 3255
rect 2290 3050 2305 3255
rect 2555 3050 2570 3255
rect 2290 3040 2345 3050
rect 2290 3020 2315 3040
rect 2335 3020 2345 3040
rect 2290 3010 2345 3020
rect 2515 3040 2570 3050
rect 2515 3020 2525 3040
rect 2545 3020 2570 3040
rect 2515 3010 2570 3020
rect 2290 2755 2305 3010
rect 2555 2755 2570 3010
rect 2645 2755 2660 3255
rect 2740 2755 2755 3255
rect 2830 3050 2845 3255
rect 3095 3050 3110 3255
rect 2830 3040 2885 3050
rect 2830 3020 2855 3040
rect 2875 3020 2885 3040
rect 2830 3010 2885 3020
rect 3055 3040 3110 3050
rect 3055 3020 3065 3040
rect 3085 3020 3110 3040
rect 3055 3010 3110 3020
rect 2830 2755 2845 3010
rect 3095 2755 3110 3010
rect 3185 2755 3200 3255
rect 3280 2755 3295 3255
rect 3370 3050 3385 3255
rect 3370 3040 3425 3050
rect 3370 3020 3395 3040
rect 3415 3020 3425 3040
rect 3370 3010 3425 3020
rect 3370 2755 3385 3010
rect -145 2455 -130 2705
rect -185 2445 -130 2455
rect -185 2425 -175 2445
rect -155 2425 -130 2445
rect -185 2415 -130 2425
rect -145 2205 -130 2415
rect -55 2205 -40 2705
rect 40 2205 55 2705
rect 130 2465 145 2705
rect 395 2465 410 2705
rect 130 2455 185 2465
rect 130 2435 155 2455
rect 175 2435 185 2455
rect 130 2425 185 2435
rect 355 2455 410 2465
rect 355 2435 365 2455
rect 385 2435 410 2455
rect 355 2425 410 2435
rect 130 2205 145 2425
rect 395 2205 410 2425
rect 485 2205 500 2705
rect 580 2205 595 2705
rect 670 2465 685 2705
rect 935 2465 950 2705
rect 670 2455 725 2465
rect 670 2435 695 2455
rect 715 2435 725 2455
rect 670 2425 725 2435
rect 895 2455 950 2465
rect 895 2435 905 2455
rect 925 2435 950 2455
rect 895 2425 950 2435
rect 670 2205 685 2425
rect 935 2205 950 2425
rect 1025 2205 1040 2705
rect 1120 2205 1135 2705
rect 1210 2465 1225 2705
rect 1475 2465 1490 2705
rect 1210 2455 1265 2465
rect 1210 2435 1235 2455
rect 1255 2435 1265 2455
rect 1210 2425 1265 2435
rect 1435 2455 1490 2465
rect 1435 2435 1445 2455
rect 1465 2435 1490 2455
rect 1435 2425 1490 2435
rect 1210 2205 1225 2425
rect 1475 2205 1490 2425
rect 1565 2205 1580 2705
rect 1660 2205 1675 2705
rect 1750 2465 1765 2705
rect 2015 2465 2030 2705
rect 1750 2455 1805 2465
rect 1750 2435 1775 2455
rect 1795 2435 1805 2455
rect 1750 2425 1805 2435
rect 1975 2455 2030 2465
rect 1975 2435 1985 2455
rect 2005 2435 2030 2455
rect 1975 2425 2030 2435
rect 1750 2205 1765 2425
rect 2015 2205 2030 2425
rect 2105 2205 2120 2705
rect 2200 2205 2215 2705
rect 2290 2465 2305 2705
rect 2555 2465 2570 2705
rect 2290 2455 2345 2465
rect 2290 2435 2315 2455
rect 2335 2435 2345 2455
rect 2290 2425 2345 2435
rect 2515 2455 2570 2465
rect 2515 2435 2525 2455
rect 2545 2435 2570 2455
rect 2515 2425 2570 2435
rect 2290 2205 2305 2425
rect 2555 2205 2570 2425
rect 2645 2205 2660 2705
rect 2740 2205 2755 2705
rect 2830 2465 2845 2705
rect 3095 2465 3110 2705
rect 2830 2455 2885 2465
rect 2830 2435 2855 2455
rect 2875 2435 2885 2455
rect 2830 2425 2885 2435
rect 3055 2455 3110 2465
rect 3055 2435 3065 2455
rect 3085 2435 3110 2455
rect 3055 2425 3110 2435
rect 2830 2205 2845 2425
rect 3095 2205 3110 2425
rect 3185 2205 3200 2705
rect 3280 2205 3295 2705
rect 3370 2465 3385 2705
rect 3370 2455 3425 2465
rect 3370 2435 3395 2455
rect 3415 2435 3425 2455
rect 3370 2425 3425 2435
rect 3370 2205 3385 2425
rect -145 1905 -130 2155
rect -185 1895 -130 1905
rect -185 1875 -175 1895
rect -155 1875 -130 1895
rect -185 1865 -130 1875
rect -145 1655 -130 1865
rect -55 1655 -40 2155
rect 40 1655 55 2155
rect 130 1915 145 2155
rect 395 1915 410 2155
rect 130 1905 185 1915
rect 130 1885 155 1905
rect 175 1885 185 1905
rect 130 1875 185 1885
rect 355 1905 410 1915
rect 355 1885 365 1905
rect 385 1885 410 1905
rect 355 1875 410 1885
rect 130 1655 145 1875
rect 395 1655 410 1875
rect 485 1655 500 2155
rect 580 1655 595 2155
rect 670 1915 685 2155
rect 935 1915 950 2155
rect 670 1905 725 1915
rect 670 1885 695 1905
rect 715 1885 725 1905
rect 670 1875 725 1885
rect 895 1905 950 1915
rect 895 1885 905 1905
rect 925 1885 950 1905
rect 895 1875 950 1885
rect 670 1655 685 1875
rect 935 1655 950 1875
rect 1025 1655 1040 2155
rect 1120 1655 1135 2155
rect 1210 1915 1225 2155
rect 1475 1915 1490 2155
rect 1210 1905 1265 1915
rect 1210 1885 1235 1905
rect 1255 1885 1265 1905
rect 1210 1875 1265 1885
rect 1435 1905 1490 1915
rect 1435 1885 1445 1905
rect 1465 1885 1490 1905
rect 1435 1875 1490 1885
rect 1210 1655 1225 1875
rect 1475 1655 1490 1875
rect 1565 1655 1580 2155
rect 1660 1655 1675 2155
rect 1750 1915 1765 2155
rect 2015 1915 2030 2155
rect 1750 1905 1805 1915
rect 1750 1885 1775 1905
rect 1795 1885 1805 1905
rect 1750 1875 1805 1885
rect 1975 1905 2030 1915
rect 1975 1885 1985 1905
rect 2005 1885 2030 1905
rect 1975 1875 2030 1885
rect 1750 1655 1765 1875
rect 2015 1655 2030 1875
rect 2105 1655 2120 2155
rect 2200 1655 2215 2155
rect 2290 1915 2305 2155
rect 2555 1915 2570 2155
rect 2290 1905 2345 1915
rect 2290 1885 2315 1905
rect 2335 1885 2345 1905
rect 2290 1875 2345 1885
rect 2515 1905 2570 1915
rect 2515 1885 2525 1905
rect 2545 1885 2570 1905
rect 2515 1875 2570 1885
rect 2290 1655 2305 1875
rect 2555 1655 2570 1875
rect 2645 1655 2660 2155
rect 2740 1655 2755 2155
rect 2830 1915 2845 2155
rect 3095 1915 3110 2155
rect 2830 1905 2885 1915
rect 2830 1885 2855 1905
rect 2875 1885 2885 1905
rect 2830 1875 2885 1885
rect 3055 1905 3110 1915
rect 3055 1885 3065 1905
rect 3085 1885 3110 1905
rect 3055 1875 3110 1885
rect 2830 1655 2845 1875
rect 3095 1655 3110 1875
rect 3185 1655 3200 2155
rect 3280 1655 3295 2155
rect 3370 1915 3385 2155
rect 3370 1905 3425 1915
rect 3370 1885 3395 1905
rect 3415 1885 3425 1905
rect 3370 1875 3425 1885
rect 3370 1655 3385 1875
rect -145 1355 -130 1605
rect -185 1345 -130 1355
rect -185 1325 -175 1345
rect -155 1325 -130 1345
rect -185 1315 -130 1325
rect -145 1105 -130 1315
rect -55 1105 -40 1605
rect 40 1105 55 1605
rect 130 1365 145 1605
rect 395 1365 410 1605
rect 130 1355 185 1365
rect 130 1335 155 1355
rect 175 1335 185 1355
rect 130 1325 185 1335
rect 355 1355 410 1365
rect 355 1335 365 1355
rect 385 1335 410 1355
rect 355 1325 410 1335
rect 130 1105 145 1325
rect 395 1105 410 1325
rect 485 1105 500 1605
rect 580 1105 595 1605
rect 670 1365 685 1605
rect 935 1365 950 1605
rect 670 1355 725 1365
rect 670 1335 695 1355
rect 715 1335 725 1355
rect 670 1325 725 1335
rect 895 1355 950 1365
rect 895 1335 905 1355
rect 925 1335 950 1355
rect 895 1325 950 1335
rect 670 1105 685 1325
rect 935 1105 950 1325
rect 1025 1105 1040 1605
rect 1120 1105 1135 1605
rect 1210 1365 1225 1605
rect 1475 1365 1490 1605
rect 1210 1355 1265 1365
rect 1210 1335 1235 1355
rect 1255 1335 1265 1355
rect 1210 1325 1265 1335
rect 1435 1355 1490 1365
rect 1435 1335 1445 1355
rect 1465 1335 1490 1355
rect 1435 1325 1490 1335
rect 1210 1105 1225 1325
rect 1475 1105 1490 1325
rect 1565 1105 1580 1605
rect 1660 1105 1675 1605
rect 1750 1365 1765 1605
rect 2015 1365 2030 1605
rect 1750 1355 1805 1365
rect 1750 1335 1775 1355
rect 1795 1335 1805 1355
rect 1750 1325 1805 1335
rect 1975 1355 2030 1365
rect 1975 1335 1985 1355
rect 2005 1335 2030 1355
rect 1975 1325 2030 1335
rect 1750 1105 1765 1325
rect 2015 1105 2030 1325
rect 2105 1105 2120 1605
rect 2200 1105 2215 1605
rect 2290 1365 2305 1605
rect 2555 1365 2570 1605
rect 2290 1355 2345 1365
rect 2290 1335 2315 1355
rect 2335 1335 2345 1355
rect 2290 1325 2345 1335
rect 2515 1355 2570 1365
rect 2515 1335 2525 1355
rect 2545 1335 2570 1355
rect 2515 1325 2570 1335
rect 2290 1105 2305 1325
rect 2555 1105 2570 1325
rect 2645 1105 2660 1605
rect 2740 1105 2755 1605
rect 2830 1365 2845 1605
rect 3095 1365 3110 1605
rect 2830 1355 2885 1365
rect 2830 1335 2855 1355
rect 2875 1335 2885 1355
rect 2830 1325 2885 1335
rect 3055 1355 3110 1365
rect 3055 1335 3065 1355
rect 3085 1335 3110 1355
rect 3055 1325 3110 1335
rect 2830 1105 2845 1325
rect 3095 1105 3110 1325
rect 3185 1105 3200 1605
rect 3280 1105 3295 1605
rect 3370 1365 3385 1605
rect 3370 1355 3425 1365
rect 3370 1335 3395 1355
rect 3415 1335 3425 1355
rect 3370 1325 3425 1335
rect 3370 1105 3385 1325
rect -145 805 -130 1055
rect -185 795 -130 805
rect -185 775 -175 795
rect -155 775 -130 795
rect -185 765 -130 775
rect -145 555 -130 765
rect -55 555 -40 1055
rect 40 555 55 1055
rect 130 815 145 1055
rect 395 815 410 1055
rect 130 805 185 815
rect 130 785 155 805
rect 175 785 185 805
rect 130 775 185 785
rect 355 805 410 815
rect 355 785 365 805
rect 385 785 410 805
rect 355 775 410 785
rect 130 555 145 775
rect 395 555 410 775
rect 485 555 500 1055
rect 580 555 595 1055
rect 670 815 685 1055
rect 935 815 950 1055
rect 670 805 725 815
rect 670 785 695 805
rect 715 785 725 805
rect 670 775 725 785
rect 895 805 950 815
rect 895 785 905 805
rect 925 785 950 805
rect 895 775 950 785
rect 670 555 685 775
rect 935 555 950 775
rect 1025 555 1040 1055
rect 1120 555 1135 1055
rect 1210 815 1225 1055
rect 1475 815 1490 1055
rect 1210 805 1265 815
rect 1210 785 1235 805
rect 1255 785 1265 805
rect 1210 775 1265 785
rect 1435 805 1490 815
rect 1435 785 1445 805
rect 1465 785 1490 805
rect 1435 775 1490 785
rect 1210 555 1225 775
rect 1475 555 1490 775
rect 1565 555 1580 1055
rect 1660 555 1675 1055
rect 1750 815 1765 1055
rect 2015 815 2030 1055
rect 1750 805 1805 815
rect 1750 785 1775 805
rect 1795 785 1805 805
rect 1750 775 1805 785
rect 1975 805 2030 815
rect 1975 785 1985 805
rect 2005 785 2030 805
rect 1975 775 2030 785
rect 1750 555 1765 775
rect 2015 555 2030 775
rect 2105 555 2120 1055
rect 2200 555 2215 1055
rect 2290 815 2305 1055
rect 2555 815 2570 1055
rect 2290 805 2345 815
rect 2290 785 2315 805
rect 2335 785 2345 805
rect 2290 775 2345 785
rect 2515 805 2570 815
rect 2515 785 2525 805
rect 2545 785 2570 805
rect 2515 775 2570 785
rect 2290 555 2305 775
rect 2555 555 2570 775
rect 2645 555 2660 1055
rect 2740 555 2755 1055
rect 2830 815 2845 1055
rect 3095 815 3110 1055
rect 2830 805 2885 815
rect 2830 785 2855 805
rect 2875 785 2885 805
rect 2830 775 2885 785
rect 3055 805 3110 815
rect 3055 785 3065 805
rect 3085 785 3110 805
rect 3055 775 3110 785
rect 2830 555 2845 775
rect 3095 555 3110 775
rect 3185 555 3200 1055
rect 3280 555 3295 1055
rect 3370 815 3385 1055
rect 3370 805 3425 815
rect 3370 785 3395 805
rect 3415 785 3425 805
rect 3370 775 3425 785
rect 3370 555 3385 775
rect -145 130 -130 375
rect -185 120 -130 130
rect -185 100 -175 120
rect -155 100 -130 120
rect -185 90 -130 100
rect -145 -125 -130 90
rect -55 -125 -40 375
rect 40 -125 55 375
rect 130 130 145 375
rect 395 130 410 375
rect 130 120 185 130
rect 130 100 155 120
rect 175 100 185 120
rect 130 90 185 100
rect 355 120 410 130
rect 355 100 365 120
rect 385 100 410 120
rect 355 90 410 100
rect 130 -125 145 90
rect 395 -125 410 90
rect 485 -125 500 375
rect 580 -125 595 375
rect 670 130 685 375
rect 935 130 950 375
rect 670 120 725 130
rect 670 100 695 120
rect 715 100 725 120
rect 670 90 725 100
rect 895 120 950 130
rect 895 100 905 120
rect 925 100 950 120
rect 895 90 950 100
rect 670 -125 685 90
rect 935 -125 950 90
rect 1025 -125 1040 375
rect 1120 -125 1135 375
rect 1210 130 1225 375
rect 1475 130 1490 375
rect 1210 120 1265 130
rect 1210 100 1235 120
rect 1255 100 1265 120
rect 1210 90 1265 100
rect 1435 120 1490 130
rect 1435 100 1445 120
rect 1465 100 1490 120
rect 1435 90 1490 100
rect 1210 -125 1225 90
rect 1475 -125 1490 90
rect 1565 -125 1580 375
rect 1660 -125 1675 375
rect 1750 130 1765 375
rect 2015 130 2030 375
rect 1750 120 1805 130
rect 1750 100 1775 120
rect 1795 100 1805 120
rect 1750 90 1805 100
rect 1975 120 2030 130
rect 1975 100 1985 120
rect 2005 100 2030 120
rect 1975 90 2030 100
rect 1750 -125 1765 90
rect 2015 -125 2030 90
rect 2105 -125 2120 375
rect 2200 -125 2215 375
rect 2290 130 2305 375
rect 2555 130 2570 375
rect 2290 120 2345 130
rect 2290 100 2315 120
rect 2335 100 2345 120
rect 2290 90 2345 100
rect 2515 120 2570 130
rect 2515 100 2525 120
rect 2545 100 2570 120
rect 2515 90 2570 100
rect 2290 -125 2305 90
rect 2555 -125 2570 90
rect 2645 -125 2660 375
rect 2740 -125 2755 375
rect 2830 130 2845 375
rect 3095 130 3110 375
rect 2830 120 2885 130
rect 2830 100 2855 120
rect 2875 100 2885 120
rect 2830 90 2885 100
rect 3055 120 3110 130
rect 3055 100 3065 120
rect 3085 100 3110 120
rect 3055 90 3110 100
rect 2830 -125 2845 90
rect 3095 -125 3110 90
rect 3185 -125 3200 375
rect 3280 -125 3295 375
rect 3370 130 3385 375
rect 3370 120 3425 130
rect 3370 100 3395 120
rect 3415 100 3425 120
rect 3370 90 3425 100
rect 3370 -125 3385 90
rect 3635 -125 3650 375
rect 3725 130 3740 375
rect 3725 120 3780 130
rect 3725 100 3750 120
rect 3770 100 3780 120
rect 3725 90 3780 100
rect 3725 -125 3740 90
rect -145 -420 -130 -175
rect -185 -430 -130 -420
rect -185 -450 -175 -430
rect -155 -450 -130 -430
rect -185 -460 -130 -450
rect -145 -675 -130 -460
rect -55 -675 -40 -175
rect 40 -675 55 -175
rect 130 -420 145 -175
rect 395 -420 410 -175
rect 130 -430 185 -420
rect 130 -450 155 -430
rect 175 -450 185 -430
rect 130 -460 185 -450
rect 355 -430 410 -420
rect 355 -450 365 -430
rect 385 -450 410 -430
rect 355 -460 410 -450
rect 130 -675 145 -460
rect 395 -675 410 -460
rect 485 -675 500 -175
rect 580 -675 595 -175
rect 670 -420 685 -175
rect 935 -420 950 -175
rect 670 -430 725 -420
rect 670 -450 695 -430
rect 715 -450 725 -430
rect 670 -460 725 -450
rect 895 -430 950 -420
rect 895 -450 905 -430
rect 925 -450 950 -430
rect 895 -460 950 -450
rect 670 -675 685 -460
rect 935 -675 950 -460
rect 1025 -675 1040 -175
rect 1120 -675 1135 -175
rect 1210 -420 1225 -175
rect 1475 -420 1490 -175
rect 1210 -430 1265 -420
rect 1210 -450 1235 -430
rect 1255 -450 1265 -430
rect 1210 -460 1265 -450
rect 1435 -430 1490 -420
rect 1435 -450 1445 -430
rect 1465 -450 1490 -430
rect 1435 -460 1490 -450
rect 1210 -675 1225 -460
rect 1475 -675 1490 -460
rect 1565 -675 1580 -175
rect 1660 -675 1675 -175
rect 1750 -420 1765 -175
rect 2015 -420 2030 -175
rect 1750 -430 1805 -420
rect 1750 -450 1775 -430
rect 1795 -450 1805 -430
rect 1750 -460 1805 -450
rect 1975 -430 2030 -420
rect 1975 -450 1985 -430
rect 2005 -450 2030 -430
rect 1975 -460 2030 -450
rect 1750 -675 1765 -460
rect 2015 -675 2030 -460
rect 2105 -675 2120 -175
rect 2200 -675 2215 -175
rect 2290 -420 2305 -175
rect 2555 -420 2570 -175
rect 2290 -430 2345 -420
rect 2290 -450 2315 -430
rect 2335 -450 2345 -430
rect 2290 -460 2345 -450
rect 2515 -430 2570 -420
rect 2515 -450 2525 -430
rect 2545 -450 2570 -430
rect 2515 -460 2570 -450
rect 2290 -675 2305 -460
rect 2555 -675 2570 -460
rect 2645 -675 2660 -175
rect 2740 -675 2755 -175
rect 2830 -420 2845 -175
rect 3095 -420 3110 -175
rect 2830 -430 2885 -420
rect 2830 -450 2855 -430
rect 2875 -450 2885 -430
rect 2830 -460 2885 -450
rect 3055 -430 3110 -420
rect 3055 -450 3065 -430
rect 3085 -450 3110 -430
rect 3055 -460 3110 -450
rect 2830 -675 2845 -460
rect 3095 -675 3110 -460
rect 3185 -675 3200 -175
rect 3280 -675 3295 -175
rect 3370 -420 3385 -175
rect 3370 -430 3425 -420
rect 3370 -450 3395 -430
rect 3415 -450 3425 -430
rect 3370 -460 3425 -450
rect 3370 -675 3385 -460
rect 3635 -675 3650 -175
rect 3725 -420 3740 -175
rect 3725 -430 3780 -420
rect 3725 -450 3750 -430
rect 3770 -450 3780 -430
rect 3725 -460 3780 -450
rect 3725 -675 3740 -460
rect -145 -970 -130 -725
rect -185 -980 -130 -970
rect -185 -1000 -175 -980
rect -155 -1000 -130 -980
rect -185 -1010 -130 -1000
rect -145 -1225 -130 -1010
rect -55 -1225 -40 -725
rect 40 -1225 55 -725
rect 130 -970 145 -725
rect 395 -970 410 -725
rect 130 -980 185 -970
rect 130 -1000 155 -980
rect 175 -1000 185 -980
rect 130 -1010 185 -1000
rect 355 -980 410 -970
rect 355 -1000 365 -980
rect 385 -1000 410 -980
rect 355 -1010 410 -1000
rect 130 -1225 145 -1010
rect 395 -1225 410 -1010
rect 485 -1225 500 -725
rect 580 -1225 595 -725
rect 670 -970 685 -725
rect 935 -970 950 -725
rect 670 -980 725 -970
rect 670 -1000 695 -980
rect 715 -1000 725 -980
rect 670 -1010 725 -1000
rect 895 -980 950 -970
rect 895 -1000 905 -980
rect 925 -1000 950 -980
rect 895 -1010 950 -1000
rect 670 -1225 685 -1010
rect 935 -1225 950 -1010
rect 1025 -1225 1040 -725
rect 1120 -1225 1135 -725
rect 1210 -970 1225 -725
rect 1475 -970 1490 -725
rect 1210 -980 1265 -970
rect 1210 -1000 1235 -980
rect 1255 -1000 1265 -980
rect 1210 -1010 1265 -1000
rect 1435 -980 1490 -970
rect 1435 -1000 1445 -980
rect 1465 -1000 1490 -980
rect 1435 -1010 1490 -1000
rect 1210 -1225 1225 -1010
rect 1475 -1225 1490 -1010
rect 1565 -1225 1580 -725
rect 1660 -1225 1675 -725
rect 1750 -970 1765 -725
rect 2015 -970 2030 -725
rect 1750 -980 1805 -970
rect 1750 -1000 1775 -980
rect 1795 -1000 1805 -980
rect 1750 -1010 1805 -1000
rect 1975 -980 2030 -970
rect 1975 -1000 1985 -980
rect 2005 -1000 2030 -980
rect 1975 -1010 2030 -1000
rect 1750 -1225 1765 -1010
rect 2015 -1225 2030 -1010
rect 2105 -1225 2120 -725
rect 2200 -1225 2215 -725
rect 2290 -970 2305 -725
rect 2555 -970 2570 -725
rect 2290 -980 2345 -970
rect 2290 -1000 2315 -980
rect 2335 -1000 2345 -980
rect 2290 -1010 2345 -1000
rect 2515 -980 2570 -970
rect 2515 -1000 2525 -980
rect 2545 -1000 2570 -980
rect 2515 -1010 2570 -1000
rect 2290 -1225 2305 -1010
rect 2555 -1225 2570 -1010
rect 2645 -1225 2660 -725
rect 2740 -1225 2755 -725
rect 2830 -970 2845 -725
rect 3095 -970 3110 -725
rect 2830 -980 2885 -970
rect 2830 -1000 2855 -980
rect 2875 -1000 2885 -980
rect 2830 -1010 2885 -1000
rect 3055 -980 3110 -970
rect 3055 -1000 3065 -980
rect 3085 -1000 3110 -980
rect 3055 -1010 3110 -1000
rect 2830 -1225 2845 -1010
rect 3095 -1225 3110 -1010
rect 3185 -1225 3200 -725
rect 3280 -1225 3295 -725
rect 3370 -970 3385 -725
rect 3370 -980 3425 -970
rect 3370 -1000 3395 -980
rect 3415 -1000 3425 -980
rect 3370 -1010 3425 -1000
rect 3370 -1225 3385 -1010
rect 3635 -1225 3650 -725
rect 3725 -970 3740 -725
rect 3725 -980 3780 -970
rect 3725 -1000 3750 -980
rect 3770 -1000 3780 -980
rect 3725 -1010 3780 -1000
rect 3725 -1225 3740 -1010
rect -145 -1520 -130 -1275
rect -185 -1530 -130 -1520
rect -185 -1550 -175 -1530
rect -155 -1550 -130 -1530
rect -185 -1560 -130 -1550
rect -145 -1775 -130 -1560
rect -55 -1775 -40 -1275
rect 40 -1775 55 -1275
rect 130 -1520 145 -1275
rect 395 -1520 410 -1275
rect 130 -1530 185 -1520
rect 130 -1550 155 -1530
rect 175 -1550 185 -1530
rect 130 -1560 185 -1550
rect 355 -1530 410 -1520
rect 355 -1550 365 -1530
rect 385 -1550 410 -1530
rect 355 -1560 410 -1550
rect 130 -1775 145 -1560
rect 395 -1775 410 -1560
rect 485 -1775 500 -1275
rect 580 -1775 595 -1275
rect 670 -1520 685 -1275
rect 935 -1520 950 -1275
rect 670 -1530 725 -1520
rect 670 -1550 695 -1530
rect 715 -1550 725 -1530
rect 670 -1560 725 -1550
rect 895 -1530 950 -1520
rect 895 -1550 905 -1530
rect 925 -1550 950 -1530
rect 895 -1560 950 -1550
rect 670 -1775 685 -1560
rect 935 -1775 950 -1560
rect 1025 -1775 1040 -1275
rect 1120 -1775 1135 -1275
rect 1210 -1520 1225 -1275
rect 1475 -1520 1490 -1275
rect 1210 -1530 1265 -1520
rect 1210 -1550 1235 -1530
rect 1255 -1550 1265 -1530
rect 1210 -1560 1265 -1550
rect 1435 -1530 1490 -1520
rect 1435 -1550 1445 -1530
rect 1465 -1550 1490 -1530
rect 1435 -1560 1490 -1550
rect 1210 -1775 1225 -1560
rect 1475 -1775 1490 -1560
rect 1565 -1775 1580 -1275
rect 1660 -1775 1675 -1275
rect 1750 -1520 1765 -1275
rect 2015 -1520 2030 -1275
rect 1750 -1530 1805 -1520
rect 1750 -1550 1775 -1530
rect 1795 -1550 1805 -1530
rect 1750 -1560 1805 -1550
rect 1975 -1530 2030 -1520
rect 1975 -1550 1985 -1530
rect 2005 -1550 2030 -1530
rect 1975 -1560 2030 -1550
rect 1750 -1775 1765 -1560
rect 2015 -1775 2030 -1560
rect 2105 -1775 2120 -1275
rect 2200 -1775 2215 -1275
rect 2290 -1520 2305 -1275
rect 2555 -1520 2570 -1275
rect 2290 -1530 2345 -1520
rect 2290 -1550 2315 -1530
rect 2335 -1550 2345 -1530
rect 2290 -1560 2345 -1550
rect 2515 -1530 2570 -1520
rect 2515 -1550 2525 -1530
rect 2545 -1550 2570 -1530
rect 2515 -1560 2570 -1550
rect 2290 -1775 2305 -1560
rect 2555 -1775 2570 -1560
rect 2645 -1775 2660 -1275
rect 2740 -1775 2755 -1275
rect 2830 -1520 2845 -1275
rect 3095 -1520 3110 -1275
rect 2830 -1530 2885 -1520
rect 2830 -1550 2855 -1530
rect 2875 -1550 2885 -1530
rect 2830 -1560 2885 -1550
rect 3055 -1530 3110 -1520
rect 3055 -1550 3065 -1530
rect 3085 -1550 3110 -1530
rect 3055 -1560 3110 -1550
rect 2830 -1775 2845 -1560
rect 3095 -1775 3110 -1560
rect 3185 -1775 3200 -1275
rect 3280 -1775 3295 -1275
rect 3370 -1520 3385 -1275
rect 3370 -1530 3425 -1520
rect 3370 -1550 3395 -1530
rect 3415 -1550 3425 -1530
rect 3370 -1560 3425 -1550
rect 3370 -1775 3385 -1560
rect 3635 -1775 3650 -1275
rect 3725 -1520 3740 -1275
rect 3725 -1530 3780 -1520
rect 3725 -1550 3750 -1530
rect 3770 -1550 3780 -1530
rect 3725 -1560 3780 -1550
rect 3725 -1775 3740 -1560
rect -145 -2050 -130 -1825
rect -185 -2060 -130 -2050
rect -185 -2080 -175 -2060
rect -155 -2080 -130 -2060
rect -185 -2090 -130 -2080
rect -145 -2325 -130 -2090
rect -55 -2325 -40 -1825
rect 40 -2325 55 -1825
rect 130 -2050 145 -1825
rect 130 -2060 185 -2050
rect 130 -2080 155 -2060
rect 175 -2080 185 -2060
rect 130 -2090 185 -2080
rect 130 -2325 145 -2090
rect 395 -2325 410 -1825
rect 485 -2050 500 -1825
rect 485 -2060 540 -2050
rect 485 -2080 510 -2060
rect 530 -2080 540 -2060
rect 485 -2090 540 -2080
rect 485 -2325 500 -2090
rect 580 -2325 595 -1825
rect 670 -2050 685 -1825
rect 670 -2060 725 -2050
rect 670 -2080 695 -2060
rect 715 -2080 725 -2060
rect 670 -2090 725 -2080
rect 670 -2325 685 -2090
rect 935 -2325 950 -1825
rect 1025 -2050 1040 -1825
rect 1025 -2060 1080 -2050
rect 1025 -2080 1050 -2060
rect 1070 -2080 1080 -2060
rect 1025 -2090 1080 -2080
rect 1025 -2325 1040 -2090
rect 1120 -2325 1135 -1825
rect 1210 -2050 1225 -1825
rect 1210 -2060 1265 -2050
rect 1210 -2080 1235 -2060
rect 1255 -2080 1265 -2060
rect 1210 -2090 1265 -2080
rect 1210 -2325 1225 -2090
rect 1475 -2325 1490 -1825
rect 1565 -2050 1580 -1825
rect 1565 -2060 1620 -2050
rect 1565 -2080 1590 -2060
rect 1610 -2080 1620 -2060
rect 1565 -2090 1620 -2080
rect 1565 -2325 1580 -2090
rect 1660 -2325 1675 -1825
rect 1750 -2050 1765 -1825
rect 1750 -2060 1805 -2050
rect 1750 -2080 1775 -2060
rect 1795 -2080 1805 -2060
rect 1750 -2090 1805 -2080
rect 1750 -2325 1765 -2090
rect 2015 -2325 2030 -1825
rect 2105 -2050 2120 -1825
rect 2105 -2060 2160 -2050
rect 2105 -2080 2130 -2060
rect 2150 -2080 2160 -2060
rect 2105 -2090 2160 -2080
rect 2105 -2325 2120 -2090
rect 2200 -2325 2215 -1825
rect 2290 -2050 2305 -1825
rect 2290 -2060 2345 -2050
rect 2290 -2080 2315 -2060
rect 2335 -2080 2345 -2060
rect 2290 -2090 2345 -2080
rect 2290 -2325 2305 -2090
rect 2555 -2325 2570 -1825
rect 2645 -2050 2660 -1825
rect 2645 -2060 2700 -2050
rect 2645 -2080 2670 -2060
rect 2690 -2080 2700 -2060
rect 2645 -2090 2700 -2080
rect 2645 -2325 2660 -2090
rect 2740 -2325 2755 -1825
rect 2830 -2050 2845 -1825
rect 2830 -2060 2885 -2050
rect 2830 -2080 2855 -2060
rect 2875 -2080 2885 -2060
rect 2830 -2090 2885 -2080
rect 2830 -2325 2845 -2090
rect 3095 -2325 3110 -1825
rect 3185 -2050 3200 -1825
rect 3185 -2060 3240 -2050
rect 3185 -2080 3210 -2060
rect 3230 -2080 3240 -2060
rect 3185 -2090 3240 -2080
rect 3185 -2325 3200 -2090
rect 3280 -2325 3295 -1825
rect 3370 -2050 3385 -1825
rect 3370 -2060 3425 -2050
rect 3370 -2080 3395 -2060
rect 3415 -2080 3425 -2060
rect 3370 -2090 3425 -2080
rect 3370 -2325 3385 -2090
rect 3635 -2325 3650 -1825
rect 3725 -2050 3740 -1825
rect 3725 -2060 3780 -2050
rect 3725 -2080 3750 -2060
rect 3770 -2080 3780 -2060
rect 3725 -2090 3780 -2080
rect 3725 -2325 3740 -2090
rect -145 -2665 -130 -2460
rect -185 -2675 -130 -2665
rect -185 -2695 -175 -2675
rect -155 -2695 -130 -2675
rect -185 -2705 -130 -2695
rect -145 -2960 -130 -2705
rect -55 -2960 -40 -2460
rect 40 -2960 55 -2460
rect 130 -2665 145 -2460
rect 395 -2665 410 -2460
rect 130 -2675 185 -2665
rect 130 -2695 155 -2675
rect 175 -2695 185 -2675
rect 130 -2705 185 -2695
rect 355 -2675 410 -2665
rect 355 -2695 365 -2675
rect 385 -2695 410 -2675
rect 355 -2705 410 -2695
rect 130 -2960 145 -2705
rect 395 -2960 410 -2705
rect 485 -2960 500 -2460
rect 580 -2960 595 -2460
rect 670 -2665 685 -2460
rect 935 -2665 950 -2460
rect 670 -2675 725 -2665
rect 670 -2695 695 -2675
rect 715 -2695 725 -2675
rect 670 -2705 725 -2695
rect 895 -2675 950 -2665
rect 895 -2695 905 -2675
rect 925 -2695 950 -2675
rect 895 -2705 950 -2695
rect 670 -2960 685 -2705
rect 935 -2960 950 -2705
rect 1025 -2960 1040 -2460
rect 1120 -2960 1135 -2460
rect 1210 -2665 1225 -2460
rect 1475 -2665 1490 -2460
rect 1210 -2675 1265 -2665
rect 1210 -2695 1235 -2675
rect 1255 -2695 1265 -2675
rect 1210 -2705 1265 -2695
rect 1435 -2675 1490 -2665
rect 1435 -2695 1445 -2675
rect 1465 -2695 1490 -2675
rect 1435 -2705 1490 -2695
rect 1210 -2960 1225 -2705
rect 1475 -2960 1490 -2705
rect 1565 -2960 1580 -2460
rect 1660 -2960 1675 -2460
rect 1750 -2665 1765 -2460
rect 2015 -2665 2030 -2460
rect 1750 -2675 1805 -2665
rect 1750 -2695 1775 -2675
rect 1795 -2695 1805 -2675
rect 1750 -2705 1805 -2695
rect 1975 -2675 2030 -2665
rect 1975 -2695 1985 -2675
rect 2005 -2695 2030 -2675
rect 1975 -2705 2030 -2695
rect 1750 -2960 1765 -2705
rect 2015 -2960 2030 -2705
rect 2105 -2960 2120 -2460
rect 2200 -2960 2215 -2460
rect 2290 -2665 2305 -2460
rect 2555 -2665 2570 -2460
rect 2290 -2675 2345 -2665
rect 2290 -2695 2315 -2675
rect 2335 -2695 2345 -2675
rect 2290 -2705 2345 -2695
rect 2515 -2675 2570 -2665
rect 2515 -2695 2525 -2675
rect 2545 -2695 2570 -2675
rect 2515 -2705 2570 -2695
rect 2290 -2960 2305 -2705
rect 2555 -2960 2570 -2705
rect 2645 -2960 2660 -2460
rect 2740 -2960 2755 -2460
rect 2830 -2665 2845 -2460
rect 3095 -2665 3110 -2460
rect 2830 -2675 2885 -2665
rect 2830 -2695 2855 -2675
rect 2875 -2695 2885 -2675
rect 2830 -2705 2885 -2695
rect 3055 -2675 3110 -2665
rect 3055 -2695 3065 -2675
rect 3085 -2695 3110 -2675
rect 3055 -2705 3110 -2695
rect 2830 -2960 2845 -2705
rect 3095 -2960 3110 -2705
rect 3185 -2960 3200 -2460
rect 3280 -2960 3295 -2460
rect 3370 -2665 3385 -2460
rect 3370 -2675 3425 -2665
rect 3370 -2695 3395 -2675
rect 3415 -2695 3425 -2675
rect 3370 -2705 3425 -2695
rect 3370 -2960 3385 -2705
rect 3635 -2960 3650 -2460
rect 3725 -2665 3740 -2460
rect 3725 -2675 3780 -2665
rect 3725 -2695 3750 -2675
rect 3770 -2695 3780 -2675
rect 3725 -2705 3780 -2695
rect 3725 -2960 3740 -2705
rect -145 -3260 -130 -3010
rect -185 -3270 -130 -3260
rect -185 -3290 -175 -3270
rect -155 -3290 -130 -3270
rect -185 -3300 -130 -3290
rect -145 -3510 -130 -3300
rect -55 -3510 -40 -3010
rect 40 -3510 55 -3010
rect 130 -3250 145 -3010
rect 395 -3250 410 -3010
rect 130 -3260 185 -3250
rect 130 -3280 155 -3260
rect 175 -3280 185 -3260
rect 130 -3290 185 -3280
rect 355 -3260 410 -3250
rect 355 -3280 365 -3260
rect 385 -3280 410 -3260
rect 355 -3290 410 -3280
rect 130 -3510 145 -3290
rect 395 -3510 410 -3290
rect 485 -3510 500 -3010
rect 580 -3510 595 -3010
rect 670 -3250 685 -3010
rect 935 -3250 950 -3010
rect 670 -3260 725 -3250
rect 670 -3280 695 -3260
rect 715 -3280 725 -3260
rect 670 -3290 725 -3280
rect 895 -3260 950 -3250
rect 895 -3280 905 -3260
rect 925 -3280 950 -3260
rect 895 -3290 950 -3280
rect 670 -3510 685 -3290
rect 935 -3510 950 -3290
rect 1025 -3510 1040 -3010
rect 1120 -3510 1135 -3010
rect 1210 -3250 1225 -3010
rect 1475 -3250 1490 -3010
rect 1210 -3260 1265 -3250
rect 1210 -3280 1235 -3260
rect 1255 -3280 1265 -3260
rect 1210 -3290 1265 -3280
rect 1435 -3260 1490 -3250
rect 1435 -3280 1445 -3260
rect 1465 -3280 1490 -3260
rect 1435 -3290 1490 -3280
rect 1210 -3510 1225 -3290
rect 1475 -3510 1490 -3290
rect 1565 -3510 1580 -3010
rect 1660 -3510 1675 -3010
rect 1750 -3250 1765 -3010
rect 2015 -3250 2030 -3010
rect 1750 -3260 1805 -3250
rect 1750 -3280 1775 -3260
rect 1795 -3280 1805 -3260
rect 1750 -3290 1805 -3280
rect 1975 -3260 2030 -3250
rect 1975 -3280 1985 -3260
rect 2005 -3280 2030 -3260
rect 1975 -3290 2030 -3280
rect 1750 -3510 1765 -3290
rect 2015 -3510 2030 -3290
rect 2105 -3510 2120 -3010
rect 2200 -3510 2215 -3010
rect 2290 -3250 2305 -3010
rect 2555 -3250 2570 -3010
rect 2290 -3260 2345 -3250
rect 2290 -3280 2315 -3260
rect 2335 -3280 2345 -3260
rect 2290 -3290 2345 -3280
rect 2515 -3260 2570 -3250
rect 2515 -3280 2525 -3260
rect 2545 -3280 2570 -3260
rect 2515 -3290 2570 -3280
rect 2290 -3510 2305 -3290
rect 2555 -3510 2570 -3290
rect 2645 -3510 2660 -3010
rect 2740 -3510 2755 -3010
rect 2830 -3250 2845 -3010
rect 3095 -3250 3110 -3010
rect 2830 -3260 2885 -3250
rect 2830 -3280 2855 -3260
rect 2875 -3280 2885 -3260
rect 2830 -3290 2885 -3280
rect 3055 -3260 3110 -3250
rect 3055 -3280 3065 -3260
rect 3085 -3280 3110 -3260
rect 3055 -3290 3110 -3280
rect 2830 -3510 2845 -3290
rect 3095 -3510 3110 -3290
rect 3185 -3510 3200 -3010
rect 3280 -3510 3295 -3010
rect 3370 -3250 3385 -3010
rect 3370 -3260 3425 -3250
rect 3370 -3280 3395 -3260
rect 3415 -3280 3425 -3260
rect 3370 -3290 3425 -3280
rect 3370 -3510 3385 -3290
rect 3635 -3510 3650 -3010
rect 3725 -3250 3740 -3010
rect 3725 -3260 3780 -3250
rect 3725 -3280 3750 -3260
rect 3770 -3280 3780 -3260
rect 3725 -3290 3780 -3280
rect 3725 -3510 3740 -3290
rect -145 -3810 -130 -3560
rect -185 -3820 -130 -3810
rect -185 -3840 -175 -3820
rect -155 -3840 -130 -3820
rect -185 -3850 -130 -3840
rect -145 -4060 -130 -3850
rect -55 -4060 -40 -3560
rect 40 -4060 55 -3560
rect 130 -3800 145 -3560
rect 395 -3800 410 -3560
rect 130 -3810 185 -3800
rect 130 -3830 155 -3810
rect 175 -3830 185 -3810
rect 130 -3840 185 -3830
rect 355 -3810 410 -3800
rect 355 -3830 365 -3810
rect 385 -3830 410 -3810
rect 355 -3840 410 -3830
rect 130 -4060 145 -3840
rect 395 -4060 410 -3840
rect 485 -4060 500 -3560
rect 580 -4060 595 -3560
rect 670 -3800 685 -3560
rect 935 -3800 950 -3560
rect 670 -3810 725 -3800
rect 670 -3830 695 -3810
rect 715 -3830 725 -3810
rect 670 -3840 725 -3830
rect 895 -3810 950 -3800
rect 895 -3830 905 -3810
rect 925 -3830 950 -3810
rect 895 -3840 950 -3830
rect 670 -4060 685 -3840
rect 935 -4060 950 -3840
rect 1025 -4060 1040 -3560
rect 1120 -4060 1135 -3560
rect 1210 -3800 1225 -3560
rect 1475 -3800 1490 -3560
rect 1210 -3810 1265 -3800
rect 1210 -3830 1235 -3810
rect 1255 -3830 1265 -3810
rect 1210 -3840 1265 -3830
rect 1435 -3810 1490 -3800
rect 1435 -3830 1445 -3810
rect 1465 -3830 1490 -3810
rect 1435 -3840 1490 -3830
rect 1210 -4060 1225 -3840
rect 1475 -4060 1490 -3840
rect 1565 -4060 1580 -3560
rect 1660 -4060 1675 -3560
rect 1750 -3800 1765 -3560
rect 2015 -3800 2030 -3560
rect 1750 -3810 1805 -3800
rect 1750 -3830 1775 -3810
rect 1795 -3830 1805 -3810
rect 1750 -3840 1805 -3830
rect 1975 -3810 2030 -3800
rect 1975 -3830 1985 -3810
rect 2005 -3830 2030 -3810
rect 1975 -3840 2030 -3830
rect 1750 -4060 1765 -3840
rect 2015 -4060 2030 -3840
rect 2105 -4060 2120 -3560
rect 2200 -4060 2215 -3560
rect 2290 -3800 2305 -3560
rect 2555 -3800 2570 -3560
rect 2290 -3810 2345 -3800
rect 2290 -3830 2315 -3810
rect 2335 -3830 2345 -3810
rect 2290 -3840 2345 -3830
rect 2515 -3810 2570 -3800
rect 2515 -3830 2525 -3810
rect 2545 -3830 2570 -3810
rect 2515 -3840 2570 -3830
rect 2290 -4060 2305 -3840
rect 2555 -4060 2570 -3840
rect 2645 -4060 2660 -3560
rect 2740 -4060 2755 -3560
rect 2830 -3800 2845 -3560
rect 3095 -3800 3110 -3560
rect 2830 -3810 2885 -3800
rect 2830 -3830 2855 -3810
rect 2875 -3830 2885 -3810
rect 2830 -3840 2885 -3830
rect 3055 -3810 3110 -3800
rect 3055 -3830 3065 -3810
rect 3085 -3830 3110 -3810
rect 3055 -3840 3110 -3830
rect 2830 -4060 2845 -3840
rect 3095 -4060 3110 -3840
rect 3185 -4060 3200 -3560
rect 3280 -4060 3295 -3560
rect 3370 -3800 3385 -3560
rect 3370 -3810 3425 -3800
rect 3370 -3830 3395 -3810
rect 3415 -3830 3425 -3810
rect 3370 -3840 3425 -3830
rect 3370 -4060 3385 -3840
rect 3635 -4060 3650 -3560
rect 3725 -3800 3740 -3560
rect 3725 -3810 3780 -3800
rect 3725 -3830 3750 -3810
rect 3770 -3830 3780 -3810
rect 3725 -3840 3780 -3830
rect 3725 -4060 3740 -3840
rect -145 -4360 -130 -4110
rect -185 -4370 -130 -4360
rect -185 -4390 -175 -4370
rect -155 -4390 -130 -4370
rect -185 -4400 -130 -4390
rect -145 -4610 -130 -4400
rect -55 -4610 -40 -4110
rect 40 -4610 55 -4110
rect 130 -4350 145 -4110
rect 395 -4350 410 -4110
rect 130 -4360 185 -4350
rect 130 -4380 155 -4360
rect 175 -4380 185 -4360
rect 130 -4390 185 -4380
rect 355 -4360 410 -4350
rect 355 -4380 365 -4360
rect 385 -4380 410 -4360
rect 355 -4390 410 -4380
rect 130 -4610 145 -4390
rect 395 -4610 410 -4390
rect 485 -4610 500 -4110
rect 580 -4610 595 -4110
rect 670 -4350 685 -4110
rect 935 -4350 950 -4110
rect 670 -4360 725 -4350
rect 670 -4380 695 -4360
rect 715 -4380 725 -4360
rect 670 -4390 725 -4380
rect 895 -4360 950 -4350
rect 895 -4380 905 -4360
rect 925 -4380 950 -4360
rect 895 -4390 950 -4380
rect 670 -4610 685 -4390
rect 935 -4610 950 -4390
rect 1025 -4610 1040 -4110
rect 1120 -4610 1135 -4110
rect 1210 -4350 1225 -4110
rect 1475 -4350 1490 -4110
rect 1210 -4360 1265 -4350
rect 1210 -4380 1235 -4360
rect 1255 -4380 1265 -4360
rect 1210 -4390 1265 -4380
rect 1435 -4360 1490 -4350
rect 1435 -4380 1445 -4360
rect 1465 -4380 1490 -4360
rect 1435 -4390 1490 -4380
rect 1210 -4610 1225 -4390
rect 1475 -4610 1490 -4390
rect 1565 -4610 1580 -4110
rect 1660 -4610 1675 -4110
rect 1750 -4350 1765 -4110
rect 2015 -4350 2030 -4110
rect 1750 -4360 1805 -4350
rect 1750 -4380 1775 -4360
rect 1795 -4380 1805 -4360
rect 1750 -4390 1805 -4380
rect 1975 -4360 2030 -4350
rect 1975 -4380 1985 -4360
rect 2005 -4380 2030 -4360
rect 1975 -4390 2030 -4380
rect 1750 -4610 1765 -4390
rect 2015 -4610 2030 -4390
rect 2105 -4610 2120 -4110
rect 2200 -4610 2215 -4110
rect 2290 -4350 2305 -4110
rect 2555 -4350 2570 -4110
rect 2290 -4360 2345 -4350
rect 2290 -4380 2315 -4360
rect 2335 -4380 2345 -4360
rect 2290 -4390 2345 -4380
rect 2515 -4360 2570 -4350
rect 2515 -4380 2525 -4360
rect 2545 -4380 2570 -4360
rect 2515 -4390 2570 -4380
rect 2290 -4610 2305 -4390
rect 2555 -4610 2570 -4390
rect 2645 -4610 2660 -4110
rect 2740 -4610 2755 -4110
rect 2830 -4350 2845 -4110
rect 3095 -4350 3110 -4110
rect 2830 -4360 2885 -4350
rect 2830 -4380 2855 -4360
rect 2875 -4380 2885 -4360
rect 2830 -4390 2885 -4380
rect 3055 -4360 3110 -4350
rect 3055 -4380 3065 -4360
rect 3085 -4380 3110 -4360
rect 3055 -4390 3110 -4380
rect 2830 -4610 2845 -4390
rect 3095 -4610 3110 -4390
rect 3185 -4610 3200 -4110
rect 3280 -4610 3295 -4110
rect 3370 -4350 3385 -4110
rect 3370 -4360 3425 -4350
rect 3370 -4380 3395 -4360
rect 3415 -4380 3425 -4360
rect 3370 -4390 3425 -4380
rect 3370 -4610 3385 -4390
rect 3635 -4610 3650 -4110
rect 3725 -4350 3740 -4110
rect 3725 -4360 3780 -4350
rect 3725 -4380 3750 -4360
rect 3770 -4380 3780 -4360
rect 3725 -4390 3780 -4380
rect 3725 -4610 3740 -4390
rect -145 -4910 -130 -4660
rect -185 -4920 -130 -4910
rect -185 -4940 -175 -4920
rect -155 -4940 -130 -4920
rect -185 -4950 -130 -4940
rect -145 -5160 -130 -4950
rect -55 -5160 -40 -4660
rect 40 -5160 55 -4660
rect 130 -4900 145 -4660
rect 395 -4900 410 -4660
rect 130 -4910 185 -4900
rect 130 -4930 155 -4910
rect 175 -4930 185 -4910
rect 130 -4940 185 -4930
rect 355 -4910 410 -4900
rect 355 -4930 365 -4910
rect 385 -4930 410 -4910
rect 355 -4940 410 -4930
rect 130 -5160 145 -4940
rect 395 -5160 410 -4940
rect 485 -5160 500 -4660
rect 580 -5160 595 -4660
rect 670 -4900 685 -4660
rect 935 -4900 950 -4660
rect 670 -4910 725 -4900
rect 670 -4930 695 -4910
rect 715 -4930 725 -4910
rect 670 -4940 725 -4930
rect 895 -4910 950 -4900
rect 895 -4930 905 -4910
rect 925 -4930 950 -4910
rect 895 -4940 950 -4930
rect 670 -5160 685 -4940
rect 935 -5160 950 -4940
rect 1025 -5160 1040 -4660
rect 1120 -5160 1135 -4660
rect 1210 -4900 1225 -4660
rect 1475 -4900 1490 -4660
rect 1210 -4910 1265 -4900
rect 1210 -4930 1235 -4910
rect 1255 -4930 1265 -4910
rect 1210 -4940 1265 -4930
rect 1435 -4910 1490 -4900
rect 1435 -4930 1445 -4910
rect 1465 -4930 1490 -4910
rect 1435 -4940 1490 -4930
rect 1210 -5160 1225 -4940
rect 1475 -5160 1490 -4940
rect 1565 -5160 1580 -4660
rect 1660 -5160 1675 -4660
rect 1750 -4900 1765 -4660
rect 2015 -4900 2030 -4660
rect 1750 -4910 1805 -4900
rect 1750 -4930 1775 -4910
rect 1795 -4930 1805 -4910
rect 1750 -4940 1805 -4930
rect 1975 -4910 2030 -4900
rect 1975 -4930 1985 -4910
rect 2005 -4930 2030 -4910
rect 1975 -4940 2030 -4930
rect 1750 -5160 1765 -4940
rect 2015 -5160 2030 -4940
rect 2105 -5160 2120 -4660
rect 2200 -5160 2215 -4660
rect 2290 -4900 2305 -4660
rect 2555 -4900 2570 -4660
rect 2290 -4910 2345 -4900
rect 2290 -4930 2315 -4910
rect 2335 -4930 2345 -4910
rect 2290 -4940 2345 -4930
rect 2515 -4910 2570 -4900
rect 2515 -4930 2525 -4910
rect 2545 -4930 2570 -4910
rect 2515 -4940 2570 -4930
rect 2290 -5160 2305 -4940
rect 2555 -5160 2570 -4940
rect 2645 -5160 2660 -4660
rect 2740 -5160 2755 -4660
rect 2830 -4900 2845 -4660
rect 3095 -4900 3110 -4660
rect 2830 -4910 2885 -4900
rect 2830 -4930 2855 -4910
rect 2875 -4930 2885 -4910
rect 2830 -4940 2885 -4930
rect 3055 -4910 3110 -4900
rect 3055 -4930 3065 -4910
rect 3085 -4930 3110 -4910
rect 3055 -4940 3110 -4930
rect 2830 -5160 2845 -4940
rect 3095 -5160 3110 -4940
rect 3185 -5160 3200 -4660
rect 3280 -5160 3295 -4660
rect 3370 -4900 3385 -4660
rect 3370 -4910 3425 -4900
rect 3370 -4930 3395 -4910
rect 3415 -4930 3425 -4910
rect 3370 -4940 3425 -4930
rect 3370 -5160 3385 -4940
rect 3635 -5160 3650 -4660
rect 3725 -4900 3740 -4660
rect 3725 -4910 3780 -4900
rect 3725 -4930 3750 -4910
rect 3770 -4930 3780 -4910
rect 3725 -4940 3780 -4930
rect 3725 -5160 3740 -4940
rect -145 -5610 -130 -5365
rect -185 -5620 -130 -5610
rect -185 -5640 -175 -5620
rect -155 -5640 -130 -5620
rect -185 -5650 -130 -5640
rect -145 -5865 -130 -5650
rect -55 -5865 -40 -5365
rect 40 -5865 55 -5365
rect 130 -5610 145 -5365
rect 395 -5610 410 -5365
rect 130 -5620 185 -5610
rect 130 -5640 155 -5620
rect 175 -5640 185 -5620
rect 130 -5650 185 -5640
rect 355 -5620 410 -5610
rect 355 -5640 365 -5620
rect 385 -5640 410 -5620
rect 355 -5650 410 -5640
rect 130 -5865 145 -5650
rect 395 -5865 410 -5650
rect 485 -5865 500 -5365
rect 580 -5865 595 -5365
rect 670 -5610 685 -5365
rect 935 -5610 950 -5365
rect 670 -5620 725 -5610
rect 670 -5640 695 -5620
rect 715 -5640 725 -5620
rect 670 -5650 725 -5640
rect 895 -5620 950 -5610
rect 895 -5640 905 -5620
rect 925 -5640 950 -5620
rect 895 -5650 950 -5640
rect 670 -5865 685 -5650
rect 935 -5865 950 -5650
rect 1025 -5865 1040 -5365
rect 1120 -5865 1135 -5365
rect 1210 -5610 1225 -5365
rect 1475 -5610 1490 -5365
rect 1210 -5620 1265 -5610
rect 1210 -5640 1235 -5620
rect 1255 -5640 1265 -5620
rect 1210 -5650 1265 -5640
rect 1435 -5620 1490 -5610
rect 1435 -5640 1445 -5620
rect 1465 -5640 1490 -5620
rect 1435 -5650 1490 -5640
rect 1210 -5865 1225 -5650
rect 1475 -5865 1490 -5650
rect 1565 -5865 1580 -5365
rect 1660 -5865 1675 -5365
rect 1750 -5610 1765 -5365
rect 2015 -5610 2030 -5365
rect 1750 -5620 1805 -5610
rect 1750 -5640 1775 -5620
rect 1795 -5640 1805 -5620
rect 1750 -5650 1805 -5640
rect 1975 -5620 2030 -5610
rect 1975 -5640 1985 -5620
rect 2005 -5640 2030 -5620
rect 1975 -5650 2030 -5640
rect 1750 -5865 1765 -5650
rect 2015 -5865 2030 -5650
rect 2105 -5865 2120 -5365
rect 2200 -5865 2215 -5365
rect 2290 -5610 2305 -5365
rect 2555 -5610 2570 -5365
rect 2290 -5620 2345 -5610
rect 2290 -5640 2315 -5620
rect 2335 -5640 2345 -5620
rect 2290 -5650 2345 -5640
rect 2515 -5620 2570 -5610
rect 2515 -5640 2525 -5620
rect 2545 -5640 2570 -5620
rect 2515 -5650 2570 -5640
rect 2290 -5865 2305 -5650
rect 2555 -5865 2570 -5650
rect 2645 -5865 2660 -5365
rect 2740 -5865 2755 -5365
rect 2830 -5610 2845 -5365
rect 3095 -5610 3110 -5365
rect 2830 -5620 2885 -5610
rect 2830 -5640 2855 -5620
rect 2875 -5640 2885 -5620
rect 2830 -5650 2885 -5640
rect 3055 -5620 3110 -5610
rect 3055 -5640 3065 -5620
rect 3085 -5640 3110 -5620
rect 3055 -5650 3110 -5640
rect 2830 -5865 2845 -5650
rect 3095 -5865 3110 -5650
rect 3185 -5865 3200 -5365
rect 3280 -5865 3295 -5365
rect 3370 -5610 3385 -5365
rect 3370 -5620 3425 -5610
rect 3370 -5640 3395 -5620
rect 3415 -5640 3425 -5620
rect 3370 -5650 3425 -5640
rect 3370 -5865 3385 -5650
rect -145 -6160 -130 -5915
rect -185 -6170 -130 -6160
rect -185 -6190 -175 -6170
rect -155 -6190 -130 -6170
rect -185 -6200 -130 -6190
rect -145 -6415 -130 -6200
rect -55 -6415 -40 -5915
rect 40 -6415 55 -5915
rect 130 -6160 145 -5915
rect 395 -6160 410 -5915
rect 130 -6170 185 -6160
rect 130 -6190 155 -6170
rect 175 -6190 185 -6170
rect 130 -6200 185 -6190
rect 355 -6170 410 -6160
rect 355 -6190 365 -6170
rect 385 -6190 410 -6170
rect 355 -6200 410 -6190
rect 130 -6415 145 -6200
rect 395 -6415 410 -6200
rect 485 -6415 500 -5915
rect 580 -6415 595 -5915
rect 670 -6160 685 -5915
rect 935 -6160 950 -5915
rect 670 -6170 725 -6160
rect 670 -6190 695 -6170
rect 715 -6190 725 -6170
rect 670 -6200 725 -6190
rect 895 -6170 950 -6160
rect 895 -6190 905 -6170
rect 925 -6190 950 -6170
rect 895 -6200 950 -6190
rect 670 -6415 685 -6200
rect 935 -6415 950 -6200
rect 1025 -6415 1040 -5915
rect 1120 -6415 1135 -5915
rect 1210 -6160 1225 -5915
rect 1475 -6160 1490 -5915
rect 1210 -6170 1265 -6160
rect 1210 -6190 1235 -6170
rect 1255 -6190 1265 -6170
rect 1210 -6200 1265 -6190
rect 1435 -6170 1490 -6160
rect 1435 -6190 1445 -6170
rect 1465 -6190 1490 -6170
rect 1435 -6200 1490 -6190
rect 1210 -6415 1225 -6200
rect 1475 -6415 1490 -6200
rect 1565 -6415 1580 -5915
rect 1660 -6415 1675 -5915
rect 1750 -6160 1765 -5915
rect 2015 -6160 2030 -5915
rect 1750 -6170 1805 -6160
rect 1750 -6190 1775 -6170
rect 1795 -6190 1805 -6170
rect 1750 -6200 1805 -6190
rect 1975 -6170 2030 -6160
rect 1975 -6190 1985 -6170
rect 2005 -6190 2030 -6170
rect 1975 -6200 2030 -6190
rect 1750 -6415 1765 -6200
rect 2015 -6415 2030 -6200
rect 2105 -6415 2120 -5915
rect 2200 -6415 2215 -5915
rect 2290 -6160 2305 -5915
rect 2555 -6160 2570 -5915
rect 2290 -6170 2345 -6160
rect 2290 -6190 2315 -6170
rect 2335 -6190 2345 -6170
rect 2290 -6200 2345 -6190
rect 2515 -6170 2570 -6160
rect 2515 -6190 2525 -6170
rect 2545 -6190 2570 -6170
rect 2515 -6200 2570 -6190
rect 2290 -6415 2305 -6200
rect 2555 -6415 2570 -6200
rect 2645 -6415 2660 -5915
rect 2740 -6415 2755 -5915
rect 2830 -6160 2845 -5915
rect 3095 -6160 3110 -5915
rect 2830 -6170 2885 -6160
rect 2830 -6190 2855 -6170
rect 2875 -6190 2885 -6170
rect 2830 -6200 2885 -6190
rect 3055 -6170 3110 -6160
rect 3055 -6190 3065 -6170
rect 3085 -6190 3110 -6170
rect 3055 -6200 3110 -6190
rect 2830 -6415 2845 -6200
rect 3095 -6415 3110 -6200
rect 3185 -6415 3200 -5915
rect 3280 -6415 3295 -5915
rect 3370 -6160 3385 -5915
rect 3370 -6170 3425 -6160
rect 3370 -6190 3395 -6170
rect 3415 -6190 3425 -6170
rect 3370 -6200 3425 -6190
rect 3370 -6415 3385 -6200
rect -145 -6710 -130 -6465
rect -185 -6720 -130 -6710
rect -185 -6740 -175 -6720
rect -155 -6740 -130 -6720
rect -185 -6750 -130 -6740
rect -145 -6965 -130 -6750
rect -55 -6965 -40 -6465
rect 40 -6965 55 -6465
rect 130 -6710 145 -6465
rect 395 -6710 410 -6465
rect 130 -6720 185 -6710
rect 130 -6740 155 -6720
rect 175 -6740 185 -6720
rect 130 -6750 185 -6740
rect 355 -6720 410 -6710
rect 355 -6740 365 -6720
rect 385 -6740 410 -6720
rect 355 -6750 410 -6740
rect 130 -6965 145 -6750
rect 395 -6965 410 -6750
rect 485 -6965 500 -6465
rect 580 -6965 595 -6465
rect 670 -6710 685 -6465
rect 935 -6710 950 -6465
rect 670 -6720 725 -6710
rect 670 -6740 695 -6720
rect 715 -6740 725 -6720
rect 670 -6750 725 -6740
rect 895 -6720 950 -6710
rect 895 -6740 905 -6720
rect 925 -6740 950 -6720
rect 895 -6750 950 -6740
rect 670 -6965 685 -6750
rect 935 -6965 950 -6750
rect 1025 -6965 1040 -6465
rect 1120 -6965 1135 -6465
rect 1210 -6710 1225 -6465
rect 1475 -6710 1490 -6465
rect 1210 -6720 1265 -6710
rect 1210 -6740 1235 -6720
rect 1255 -6740 1265 -6720
rect 1210 -6750 1265 -6740
rect 1435 -6720 1490 -6710
rect 1435 -6740 1445 -6720
rect 1465 -6740 1490 -6720
rect 1435 -6750 1490 -6740
rect 1210 -6965 1225 -6750
rect 1475 -6965 1490 -6750
rect 1565 -6965 1580 -6465
rect 1660 -6965 1675 -6465
rect 1750 -6710 1765 -6465
rect 2015 -6710 2030 -6465
rect 1750 -6720 1805 -6710
rect 1750 -6740 1775 -6720
rect 1795 -6740 1805 -6720
rect 1750 -6750 1805 -6740
rect 1975 -6720 2030 -6710
rect 1975 -6740 1985 -6720
rect 2005 -6740 2030 -6720
rect 1975 -6750 2030 -6740
rect 1750 -6965 1765 -6750
rect 2015 -6965 2030 -6750
rect 2105 -6965 2120 -6465
rect 2200 -6965 2215 -6465
rect 2290 -6710 2305 -6465
rect 2555 -6710 2570 -6465
rect 2290 -6720 2345 -6710
rect 2290 -6740 2315 -6720
rect 2335 -6740 2345 -6720
rect 2290 -6750 2345 -6740
rect 2515 -6720 2570 -6710
rect 2515 -6740 2525 -6720
rect 2545 -6740 2570 -6720
rect 2515 -6750 2570 -6740
rect 2290 -6965 2305 -6750
rect 2555 -6965 2570 -6750
rect 2645 -6965 2660 -6465
rect 2740 -6965 2755 -6465
rect 2830 -6710 2845 -6465
rect 3095 -6710 3110 -6465
rect 2830 -6720 2885 -6710
rect 2830 -6740 2855 -6720
rect 2875 -6740 2885 -6720
rect 2830 -6750 2885 -6740
rect 3055 -6720 3110 -6710
rect 3055 -6740 3065 -6720
rect 3085 -6740 3110 -6720
rect 3055 -6750 3110 -6740
rect 2830 -6965 2845 -6750
rect 3095 -6965 3110 -6750
rect 3185 -6965 3200 -6465
rect 3280 -6965 3295 -6465
rect 3370 -6710 3385 -6465
rect 3370 -6720 3425 -6710
rect 3370 -6740 3395 -6720
rect 3415 -6740 3425 -6720
rect 3370 -6750 3425 -6740
rect 3370 -6965 3385 -6750
rect -145 -7260 -130 -7015
rect -185 -7270 -130 -7260
rect -185 -7290 -175 -7270
rect -155 -7290 -130 -7270
rect -185 -7300 -130 -7290
rect -145 -7515 -130 -7300
rect -55 -7515 -40 -7015
rect 40 -7515 55 -7015
rect 130 -7260 145 -7015
rect 395 -7260 410 -7015
rect 130 -7270 185 -7260
rect 130 -7290 155 -7270
rect 175 -7290 185 -7270
rect 130 -7300 185 -7290
rect 355 -7270 410 -7260
rect 355 -7290 365 -7270
rect 385 -7290 410 -7270
rect 355 -7300 410 -7290
rect 130 -7515 145 -7300
rect 395 -7515 410 -7300
rect 485 -7515 500 -7015
rect 580 -7515 595 -7015
rect 670 -7260 685 -7015
rect 935 -7260 950 -7015
rect 670 -7270 725 -7260
rect 670 -7290 695 -7270
rect 715 -7290 725 -7270
rect 670 -7300 725 -7290
rect 895 -7270 950 -7260
rect 895 -7290 905 -7270
rect 925 -7290 950 -7270
rect 895 -7300 950 -7290
rect 670 -7515 685 -7300
rect 935 -7515 950 -7300
rect 1025 -7515 1040 -7015
rect 1120 -7515 1135 -7015
rect 1210 -7260 1225 -7015
rect 1475 -7260 1490 -7015
rect 1210 -7270 1265 -7260
rect 1210 -7290 1235 -7270
rect 1255 -7290 1265 -7270
rect 1210 -7300 1265 -7290
rect 1435 -7270 1490 -7260
rect 1435 -7290 1445 -7270
rect 1465 -7290 1490 -7270
rect 1435 -7300 1490 -7290
rect 1210 -7515 1225 -7300
rect 1475 -7515 1490 -7300
rect 1565 -7515 1580 -7015
rect 1660 -7515 1675 -7015
rect 1750 -7260 1765 -7015
rect 2015 -7260 2030 -7015
rect 1750 -7270 1805 -7260
rect 1750 -7290 1775 -7270
rect 1795 -7290 1805 -7270
rect 1750 -7300 1805 -7290
rect 1975 -7270 2030 -7260
rect 1975 -7290 1985 -7270
rect 2005 -7290 2030 -7270
rect 1975 -7300 2030 -7290
rect 1750 -7515 1765 -7300
rect 2015 -7515 2030 -7300
rect 2105 -7515 2120 -7015
rect 2200 -7515 2215 -7015
rect 2290 -7260 2305 -7015
rect 2555 -7260 2570 -7015
rect 2290 -7270 2345 -7260
rect 2290 -7290 2315 -7270
rect 2335 -7290 2345 -7270
rect 2290 -7300 2345 -7290
rect 2515 -7270 2570 -7260
rect 2515 -7290 2525 -7270
rect 2545 -7290 2570 -7270
rect 2515 -7300 2570 -7290
rect 2290 -7515 2305 -7300
rect 2555 -7515 2570 -7300
rect 2645 -7515 2660 -7015
rect 2740 -7515 2755 -7015
rect 2830 -7260 2845 -7015
rect 3095 -7260 3110 -7015
rect 2830 -7270 2885 -7260
rect 2830 -7290 2855 -7270
rect 2875 -7290 2885 -7270
rect 2830 -7300 2885 -7290
rect 3055 -7270 3110 -7260
rect 3055 -7290 3065 -7270
rect 3085 -7290 3110 -7270
rect 3055 -7300 3110 -7290
rect 2830 -7515 2845 -7300
rect 3095 -7515 3110 -7300
rect 3185 -7515 3200 -7015
rect 3280 -7515 3295 -7015
rect 3370 -7260 3385 -7015
rect 3370 -7270 3425 -7260
rect 3370 -7290 3395 -7270
rect 3415 -7290 3425 -7270
rect 3370 -7300 3425 -7290
rect 3370 -7515 3385 -7300
rect -145 -8065 -130 -7565
rect -55 -7790 -40 -7565
rect -55 -7800 0 -7790
rect -55 -7820 -30 -7800
rect -10 -7820 0 -7800
rect -55 -7830 0 -7820
rect -55 -8065 -40 -7830
rect 40 -8065 55 -7565
rect 130 -7790 145 -7565
rect 130 -7800 185 -7790
rect 130 -7820 155 -7800
rect 175 -7820 185 -7800
rect 130 -7830 185 -7820
rect 130 -8065 145 -7830
rect 395 -8065 410 -7565
rect 485 -7790 500 -7565
rect 485 -7800 540 -7790
rect 485 -7820 510 -7800
rect 530 -7820 540 -7800
rect 485 -7830 540 -7820
rect 485 -8065 500 -7830
rect 580 -8065 595 -7565
rect 670 -7790 685 -7565
rect 670 -7800 725 -7790
rect 670 -7820 695 -7800
rect 715 -7820 725 -7800
rect 670 -7830 725 -7820
rect 670 -8065 685 -7830
rect 935 -8065 950 -7565
rect 1025 -7790 1040 -7565
rect 1025 -7800 1080 -7790
rect 1025 -7820 1050 -7800
rect 1070 -7820 1080 -7800
rect 1025 -7830 1080 -7820
rect 1025 -8065 1040 -7830
rect 1120 -8065 1135 -7565
rect 1210 -7790 1225 -7565
rect 1210 -7800 1265 -7790
rect 1210 -7820 1235 -7800
rect 1255 -7820 1265 -7800
rect 1210 -7830 1265 -7820
rect 1210 -8065 1225 -7830
rect 1475 -8065 1490 -7565
rect 1565 -7790 1580 -7565
rect 1565 -7800 1620 -7790
rect 1565 -7820 1590 -7800
rect 1610 -7820 1620 -7800
rect 1565 -7830 1620 -7820
rect 1565 -8065 1580 -7830
rect 1660 -8065 1675 -7565
rect 1750 -7790 1765 -7565
rect 1750 -7800 1805 -7790
rect 1750 -7820 1775 -7800
rect 1795 -7820 1805 -7800
rect 1750 -7830 1805 -7820
rect 1750 -8065 1765 -7830
rect 2015 -8065 2030 -7565
rect 2105 -7790 2120 -7565
rect 2105 -7800 2160 -7790
rect 2105 -7820 2130 -7800
rect 2150 -7820 2160 -7800
rect 2105 -7830 2160 -7820
rect 2105 -8065 2120 -7830
rect 2200 -8065 2215 -7565
rect 2290 -7790 2305 -7565
rect 2290 -7800 2345 -7790
rect 2290 -7820 2315 -7800
rect 2335 -7820 2345 -7800
rect 2290 -7830 2345 -7820
rect 2290 -8065 2305 -7830
rect 2555 -8065 2570 -7565
rect 2645 -7790 2660 -7565
rect 2645 -7800 2700 -7790
rect 2645 -7820 2670 -7800
rect 2690 -7820 2700 -7800
rect 2645 -7830 2700 -7820
rect 2645 -8065 2660 -7830
rect 2740 -8065 2755 -7565
rect 2830 -7790 2845 -7565
rect 2830 -7800 2885 -7790
rect 2830 -7820 2855 -7800
rect 2875 -7820 2885 -7800
rect 2830 -7830 2885 -7820
rect 2830 -8065 2845 -7830
rect 3095 -8065 3110 -7565
rect 3185 -7790 3200 -7565
rect 3185 -7800 3240 -7790
rect 3185 -7820 3210 -7800
rect 3230 -7820 3240 -7800
rect 3185 -7830 3240 -7820
rect 3185 -8065 3200 -7830
rect 3280 -8065 3295 -7565
rect 3370 -7790 3385 -7565
rect 3370 -7800 3425 -7790
rect 3370 -7820 3395 -7800
rect 3415 -7820 3425 -7800
rect 3370 -7830 3425 -7820
rect 3370 -8065 3385 -7830
<< polycont >>
rect -30 3020 -10 3040
rect 155 3020 175 3040
rect 365 3020 385 3040
rect 695 3020 715 3040
rect 905 3020 925 3040
rect 1235 3020 1255 3040
rect 1445 3020 1465 3040
rect 1775 3020 1795 3040
rect 1985 3020 2005 3040
rect 2315 3020 2335 3040
rect 2525 3020 2545 3040
rect 2855 3020 2875 3040
rect 3065 3020 3085 3040
rect 3395 3020 3415 3040
rect -175 2425 -155 2445
rect 155 2435 175 2455
rect 365 2435 385 2455
rect 695 2435 715 2455
rect 905 2435 925 2455
rect 1235 2435 1255 2455
rect 1445 2435 1465 2455
rect 1775 2435 1795 2455
rect 1985 2435 2005 2455
rect 2315 2435 2335 2455
rect 2525 2435 2545 2455
rect 2855 2435 2875 2455
rect 3065 2435 3085 2455
rect 3395 2435 3415 2455
rect -175 1875 -155 1895
rect 155 1885 175 1905
rect 365 1885 385 1905
rect 695 1885 715 1905
rect 905 1885 925 1905
rect 1235 1885 1255 1905
rect 1445 1885 1465 1905
rect 1775 1885 1795 1905
rect 1985 1885 2005 1905
rect 2315 1885 2335 1905
rect 2525 1885 2545 1905
rect 2855 1885 2875 1905
rect 3065 1885 3085 1905
rect 3395 1885 3415 1905
rect -175 1325 -155 1345
rect 155 1335 175 1355
rect 365 1335 385 1355
rect 695 1335 715 1355
rect 905 1335 925 1355
rect 1235 1335 1255 1355
rect 1445 1335 1465 1355
rect 1775 1335 1795 1355
rect 1985 1335 2005 1355
rect 2315 1335 2335 1355
rect 2525 1335 2545 1355
rect 2855 1335 2875 1355
rect 3065 1335 3085 1355
rect 3395 1335 3415 1355
rect -175 775 -155 795
rect 155 785 175 805
rect 365 785 385 805
rect 695 785 715 805
rect 905 785 925 805
rect 1235 785 1255 805
rect 1445 785 1465 805
rect 1775 785 1795 805
rect 1985 785 2005 805
rect 2315 785 2335 805
rect 2525 785 2545 805
rect 2855 785 2875 805
rect 3065 785 3085 805
rect 3395 785 3415 805
rect -175 100 -155 120
rect 155 100 175 120
rect 365 100 385 120
rect 695 100 715 120
rect 905 100 925 120
rect 1235 100 1255 120
rect 1445 100 1465 120
rect 1775 100 1795 120
rect 1985 100 2005 120
rect 2315 100 2335 120
rect 2525 100 2545 120
rect 2855 100 2875 120
rect 3065 100 3085 120
rect 3395 100 3415 120
rect 3750 100 3770 120
rect -175 -450 -155 -430
rect 155 -450 175 -430
rect 365 -450 385 -430
rect 695 -450 715 -430
rect 905 -450 925 -430
rect 1235 -450 1255 -430
rect 1445 -450 1465 -430
rect 1775 -450 1795 -430
rect 1985 -450 2005 -430
rect 2315 -450 2335 -430
rect 2525 -450 2545 -430
rect 2855 -450 2875 -430
rect 3065 -450 3085 -430
rect 3395 -450 3415 -430
rect 3750 -450 3770 -430
rect -175 -1000 -155 -980
rect 155 -1000 175 -980
rect 365 -1000 385 -980
rect 695 -1000 715 -980
rect 905 -1000 925 -980
rect 1235 -1000 1255 -980
rect 1445 -1000 1465 -980
rect 1775 -1000 1795 -980
rect 1985 -1000 2005 -980
rect 2315 -1000 2335 -980
rect 2525 -1000 2545 -980
rect 2855 -1000 2875 -980
rect 3065 -1000 3085 -980
rect 3395 -1000 3415 -980
rect 3750 -1000 3770 -980
rect -175 -1550 -155 -1530
rect 155 -1550 175 -1530
rect 365 -1550 385 -1530
rect 695 -1550 715 -1530
rect 905 -1550 925 -1530
rect 1235 -1550 1255 -1530
rect 1445 -1550 1465 -1530
rect 1775 -1550 1795 -1530
rect 1985 -1550 2005 -1530
rect 2315 -1550 2335 -1530
rect 2525 -1550 2545 -1530
rect 2855 -1550 2875 -1530
rect 3065 -1550 3085 -1530
rect 3395 -1550 3415 -1530
rect 3750 -1550 3770 -1530
rect -175 -2080 -155 -2060
rect 155 -2080 175 -2060
rect 510 -2080 530 -2060
rect 695 -2080 715 -2060
rect 1050 -2080 1070 -2060
rect 1235 -2080 1255 -2060
rect 1590 -2080 1610 -2060
rect 1775 -2080 1795 -2060
rect 2130 -2080 2150 -2060
rect 2315 -2080 2335 -2060
rect 2670 -2080 2690 -2060
rect 2855 -2080 2875 -2060
rect 3210 -2080 3230 -2060
rect 3395 -2080 3415 -2060
rect 3750 -2080 3770 -2060
rect -175 -2695 -155 -2675
rect 155 -2695 175 -2675
rect 365 -2695 385 -2675
rect 695 -2695 715 -2675
rect 905 -2695 925 -2675
rect 1235 -2695 1255 -2675
rect 1445 -2695 1465 -2675
rect 1775 -2695 1795 -2675
rect 1985 -2695 2005 -2675
rect 2315 -2695 2335 -2675
rect 2525 -2695 2545 -2675
rect 2855 -2695 2875 -2675
rect 3065 -2695 3085 -2675
rect 3395 -2695 3415 -2675
rect 3750 -2695 3770 -2675
rect -175 -3290 -155 -3270
rect 155 -3280 175 -3260
rect 365 -3280 385 -3260
rect 695 -3280 715 -3260
rect 905 -3280 925 -3260
rect 1235 -3280 1255 -3260
rect 1445 -3280 1465 -3260
rect 1775 -3280 1795 -3260
rect 1985 -3280 2005 -3260
rect 2315 -3280 2335 -3260
rect 2525 -3280 2545 -3260
rect 2855 -3280 2875 -3260
rect 3065 -3280 3085 -3260
rect 3395 -3280 3415 -3260
rect 3750 -3280 3770 -3260
rect -175 -3840 -155 -3820
rect 155 -3830 175 -3810
rect 365 -3830 385 -3810
rect 695 -3830 715 -3810
rect 905 -3830 925 -3810
rect 1235 -3830 1255 -3810
rect 1445 -3830 1465 -3810
rect 1775 -3830 1795 -3810
rect 1985 -3830 2005 -3810
rect 2315 -3830 2335 -3810
rect 2525 -3830 2545 -3810
rect 2855 -3830 2875 -3810
rect 3065 -3830 3085 -3810
rect 3395 -3830 3415 -3810
rect 3750 -3830 3770 -3810
rect -175 -4390 -155 -4370
rect 155 -4380 175 -4360
rect 365 -4380 385 -4360
rect 695 -4380 715 -4360
rect 905 -4380 925 -4360
rect 1235 -4380 1255 -4360
rect 1445 -4380 1465 -4360
rect 1775 -4380 1795 -4360
rect 1985 -4380 2005 -4360
rect 2315 -4380 2335 -4360
rect 2525 -4380 2545 -4360
rect 2855 -4380 2875 -4360
rect 3065 -4380 3085 -4360
rect 3395 -4380 3415 -4360
rect 3750 -4380 3770 -4360
rect -175 -4940 -155 -4920
rect 155 -4930 175 -4910
rect 365 -4930 385 -4910
rect 695 -4930 715 -4910
rect 905 -4930 925 -4910
rect 1235 -4930 1255 -4910
rect 1445 -4930 1465 -4910
rect 1775 -4930 1795 -4910
rect 1985 -4930 2005 -4910
rect 2315 -4930 2335 -4910
rect 2525 -4930 2545 -4910
rect 2855 -4930 2875 -4910
rect 3065 -4930 3085 -4910
rect 3395 -4930 3415 -4910
rect 3750 -4930 3770 -4910
rect -175 -5640 -155 -5620
rect 155 -5640 175 -5620
rect 365 -5640 385 -5620
rect 695 -5640 715 -5620
rect 905 -5640 925 -5620
rect 1235 -5640 1255 -5620
rect 1445 -5640 1465 -5620
rect 1775 -5640 1795 -5620
rect 1985 -5640 2005 -5620
rect 2315 -5640 2335 -5620
rect 2525 -5640 2545 -5620
rect 2855 -5640 2875 -5620
rect 3065 -5640 3085 -5620
rect 3395 -5640 3415 -5620
rect -175 -6190 -155 -6170
rect 155 -6190 175 -6170
rect 365 -6190 385 -6170
rect 695 -6190 715 -6170
rect 905 -6190 925 -6170
rect 1235 -6190 1255 -6170
rect 1445 -6190 1465 -6170
rect 1775 -6190 1795 -6170
rect 1985 -6190 2005 -6170
rect 2315 -6190 2335 -6170
rect 2525 -6190 2545 -6170
rect 2855 -6190 2875 -6170
rect 3065 -6190 3085 -6170
rect 3395 -6190 3415 -6170
rect -175 -6740 -155 -6720
rect 155 -6740 175 -6720
rect 365 -6740 385 -6720
rect 695 -6740 715 -6720
rect 905 -6740 925 -6720
rect 1235 -6740 1255 -6720
rect 1445 -6740 1465 -6720
rect 1775 -6740 1795 -6720
rect 1985 -6740 2005 -6720
rect 2315 -6740 2335 -6720
rect 2525 -6740 2545 -6720
rect 2855 -6740 2875 -6720
rect 3065 -6740 3085 -6720
rect 3395 -6740 3415 -6720
rect -175 -7290 -155 -7270
rect 155 -7290 175 -7270
rect 365 -7290 385 -7270
rect 695 -7290 715 -7270
rect 905 -7290 925 -7270
rect 1235 -7290 1255 -7270
rect 1445 -7290 1465 -7270
rect 1775 -7290 1795 -7270
rect 1985 -7290 2005 -7270
rect 2315 -7290 2335 -7270
rect 2525 -7290 2545 -7270
rect 2855 -7290 2875 -7270
rect 3065 -7290 3085 -7270
rect 3395 -7290 3415 -7270
rect -30 -7820 -10 -7800
rect 155 -7820 175 -7800
rect 510 -7820 530 -7800
rect 695 -7820 715 -7800
rect 1050 -7820 1070 -7800
rect 1235 -7820 1255 -7800
rect 1590 -7820 1610 -7800
rect 1775 -7820 1795 -7800
rect 2130 -7820 2150 -7800
rect 2315 -7820 2335 -7800
rect 2670 -7820 2690 -7800
rect 2855 -7820 2875 -7800
rect 3210 -7820 3230 -7800
rect 3395 -7820 3415 -7800
<< locali >>
rect -425 3785 1410 3805
rect -425 -8540 -405 3785
rect -385 3745 1320 3765
rect -385 -8500 -365 3745
rect -345 3705 870 3725
rect -345 -8460 -325 3705
rect -305 3665 780 3685
rect -305 -8420 -285 3665
rect -265 3625 330 3645
rect -265 -8380 -245 3625
rect -225 3585 240 3605
rect -225 -8340 -205 3585
rect 220 3550 240 3585
rect 310 3550 330 3625
rect 760 3550 780 3665
rect 850 3550 870 3705
rect 1300 3550 1320 3745
rect 1390 3550 1410 3785
rect 1840 3785 4020 3805
rect 1840 3550 1860 3785
rect 1930 3745 3980 3765
rect 1930 3550 1950 3745
rect 2380 3705 3940 3725
rect 2380 3550 2400 3705
rect 2470 3665 3900 3685
rect 2470 3550 2490 3665
rect 2920 3625 3860 3645
rect 2920 3550 2940 3625
rect 3010 3585 3820 3605
rect 3010 3550 3030 3585
rect 205 3540 255 3550
rect 205 3460 215 3540
rect 245 3460 255 3540
rect 205 3450 255 3460
rect 295 3540 345 3550
rect 295 3460 305 3540
rect 335 3460 345 3540
rect 295 3450 345 3460
rect 745 3540 795 3550
rect 745 3460 755 3540
rect 785 3460 795 3540
rect 745 3450 795 3460
rect 835 3540 885 3550
rect 835 3460 845 3540
rect 875 3460 885 3540
rect 835 3450 885 3460
rect 1285 3540 1335 3550
rect 1285 3460 1295 3540
rect 1325 3460 1335 3540
rect 1285 3450 1335 3460
rect 1375 3540 1425 3550
rect 1375 3460 1385 3540
rect 1415 3460 1425 3540
rect 1375 3450 1425 3460
rect 1825 3540 1875 3550
rect 1825 3460 1835 3540
rect 1865 3460 1875 3540
rect 1825 3450 1875 3460
rect 1915 3540 1965 3550
rect 1915 3460 1925 3540
rect 1955 3460 1965 3540
rect 1915 3450 1965 3460
rect 2365 3540 2415 3550
rect 2365 3460 2375 3540
rect 2405 3460 2415 3540
rect 2365 3450 2415 3460
rect 2455 3540 2505 3550
rect 2455 3460 2465 3540
rect 2495 3460 2505 3540
rect 2455 3450 2505 3460
rect 2905 3540 2955 3550
rect 2905 3460 2915 3540
rect 2945 3460 2955 3540
rect 2905 3450 2955 3460
rect 2995 3540 3045 3550
rect 2995 3460 3005 3540
rect 3035 3460 3045 3540
rect 2995 3450 3045 3460
rect -125 3290 3425 3300
rect -125 3270 -115 3290
rect -70 3280 70 3290
rect -70 3270 -60 3280
rect -125 3260 -60 3270
rect 60 3270 70 3280
rect 115 3280 425 3290
rect 115 3270 125 3280
rect 60 3260 125 3270
rect 415 3270 425 3280
rect 470 3280 610 3290
rect 470 3270 480 3280
rect 415 3260 480 3270
rect 600 3270 610 3280
rect 655 3280 965 3290
rect 655 3270 665 3280
rect 600 3260 665 3270
rect 955 3270 965 3280
rect 1010 3280 1150 3290
rect 1010 3270 1020 3280
rect 955 3260 1020 3270
rect 1140 3270 1150 3280
rect 1195 3280 1505 3290
rect 1195 3270 1205 3280
rect 1140 3260 1205 3270
rect 1495 3270 1505 3280
rect 1550 3280 1690 3290
rect 1550 3270 1560 3280
rect 1495 3260 1560 3270
rect 1680 3270 1690 3280
rect 1735 3280 2045 3290
rect 1735 3270 1745 3280
rect 1680 3260 1745 3270
rect 2035 3270 2045 3280
rect 2090 3280 2230 3290
rect 2090 3270 2100 3280
rect 2035 3260 2100 3270
rect 2220 3270 2230 3280
rect 2275 3280 2585 3290
rect 2275 3270 2285 3280
rect 2220 3260 2285 3270
rect 2575 3270 2585 3280
rect 2630 3280 2770 3290
rect 2630 3270 2640 3280
rect 2575 3260 2640 3270
rect 2760 3270 2770 3280
rect 2815 3280 3125 3290
rect 2815 3270 2825 3280
rect 2760 3260 2825 3270
rect 3115 3270 3125 3280
rect 3170 3280 3310 3290
rect 3170 3270 3180 3280
rect 3115 3260 3180 3270
rect 3300 3270 3310 3280
rect 3355 3280 3425 3290
rect 3355 3270 3365 3280
rect 3300 3260 3365 3270
rect 3405 3050 3425 3280
rect -40 3040 3425 3050
rect -40 3020 -30 3040
rect -10 3030 155 3040
rect -10 3020 0 3030
rect -40 3010 0 3020
rect 145 3020 155 3030
rect 175 3030 365 3040
rect 175 3020 185 3030
rect 145 3010 185 3020
rect 355 3020 365 3030
rect 385 3030 695 3040
rect 385 3020 395 3030
rect 355 3010 395 3020
rect 685 3020 695 3030
rect 715 3030 905 3040
rect 715 3020 725 3030
rect 685 3010 725 3020
rect 895 3020 905 3030
rect 925 3030 1235 3040
rect 925 3020 935 3030
rect 895 3010 935 3020
rect 1225 3020 1235 3030
rect 1255 3030 1445 3040
rect 1255 3020 1265 3030
rect 1225 3010 1265 3020
rect 1435 3020 1445 3030
rect 1465 3030 1775 3040
rect 1465 3020 1475 3030
rect 1435 3010 1475 3020
rect 1765 3020 1775 3030
rect 1795 3030 1985 3040
rect 1795 3020 1805 3030
rect 1765 3010 1805 3020
rect 1975 3020 1985 3030
rect 2005 3030 2315 3040
rect 2005 3020 2015 3030
rect 1975 3010 2015 3020
rect 2305 3020 2315 3030
rect 2335 3030 2525 3040
rect 2335 3020 2345 3030
rect 2305 3010 2345 3020
rect 2515 3020 2525 3030
rect 2545 3030 2855 3040
rect 2545 3020 2555 3030
rect 2515 3010 2555 3020
rect 2845 3020 2855 3030
rect 2875 3030 3065 3040
rect 2875 3020 2885 3030
rect 2845 3010 2885 3020
rect 3055 3020 3065 3030
rect 3085 3030 3395 3040
rect 3085 3020 3095 3030
rect 3055 3010 3095 3020
rect 3385 3020 3395 3030
rect 3415 3020 3425 3040
rect 3385 3010 3425 3020
rect -125 2740 -60 2750
rect -125 2720 -115 2740
rect -70 2720 -60 2740
rect -125 2710 -60 2720
rect 60 2740 125 2750
rect 60 2720 70 2740
rect 115 2720 125 2740
rect 60 2710 125 2720
rect 415 2740 480 2750
rect 415 2720 425 2740
rect 470 2720 480 2740
rect 415 2710 480 2720
rect 600 2740 665 2750
rect 600 2720 610 2740
rect 655 2720 665 2740
rect 600 2710 665 2720
rect 955 2740 1020 2750
rect 955 2720 965 2740
rect 1010 2720 1020 2740
rect 955 2710 1020 2720
rect 1140 2740 1205 2750
rect 1140 2720 1150 2740
rect 1195 2720 1205 2740
rect 1140 2710 1205 2720
rect 1495 2740 1560 2750
rect 1495 2720 1505 2740
rect 1550 2720 1560 2740
rect 1495 2710 1560 2720
rect 1680 2740 1745 2750
rect 1680 2720 1690 2740
rect 1735 2720 1745 2740
rect 1680 2710 1745 2720
rect 2035 2740 2100 2750
rect 2035 2720 2045 2740
rect 2090 2720 2100 2740
rect 2035 2710 2100 2720
rect 2220 2740 2285 2750
rect 2220 2720 2230 2740
rect 2275 2720 2285 2740
rect 2220 2710 2285 2720
rect 2575 2740 2640 2750
rect 2575 2720 2585 2740
rect 2630 2720 2640 2740
rect 2575 2710 2640 2720
rect 2760 2740 2825 2750
rect 2760 2720 2770 2740
rect 2815 2720 2825 2740
rect 2760 2710 2825 2720
rect 3115 2740 3180 2750
rect 3115 2720 3125 2740
rect 3170 2720 3180 2740
rect 3115 2710 3180 2720
rect 3300 2740 3365 2750
rect 3300 2720 3310 2740
rect 3355 2720 3365 2740
rect 3300 2710 3365 2720
rect 145 2455 185 2465
rect -185 2445 -145 2455
rect -185 2425 -175 2445
rect -155 2425 -145 2445
rect 145 2435 155 2455
rect 175 2435 185 2455
rect 145 2425 185 2435
rect -185 2415 -145 2425
rect 165 2415 185 2425
rect 355 2455 395 2465
rect 355 2435 365 2455
rect 385 2435 395 2455
rect 355 2425 395 2435
rect 685 2455 725 2465
rect 685 2435 695 2455
rect 715 2435 725 2455
rect 685 2425 725 2435
rect -185 1905 -165 2415
rect 165 2405 260 2415
rect 165 2375 195 2405
rect 250 2375 260 2405
rect 165 2365 260 2375
rect -125 2190 -60 2200
rect -125 2170 -115 2190
rect -70 2170 -60 2190
rect -125 2160 -60 2170
rect 60 2190 125 2200
rect 60 2170 70 2190
rect 115 2170 125 2190
rect 60 2160 125 2170
rect 165 1915 185 2365
rect 355 2340 375 2425
rect 280 2330 375 2340
rect 280 2300 290 2330
rect 345 2300 375 2330
rect 280 2290 375 2300
rect 145 1905 185 1915
rect -185 1895 -145 1905
rect -185 1875 -175 1895
rect -155 1875 -145 1895
rect 145 1885 155 1905
rect 175 1885 185 1905
rect 145 1875 185 1885
rect -185 1865 -145 1875
rect -185 1355 -165 1865
rect -20 1860 20 1870
rect -20 1790 -10 1860
rect 10 1790 20 1860
rect -20 1780 20 1790
rect -125 1640 -60 1650
rect -125 1620 -115 1640
rect -70 1620 -60 1640
rect -125 1610 -60 1620
rect 60 1640 125 1650
rect 60 1620 70 1640
rect 115 1620 125 1640
rect 60 1610 125 1620
rect 165 1365 185 1875
rect 145 1355 185 1365
rect -185 1345 -145 1355
rect -185 1325 -175 1345
rect -155 1325 -145 1345
rect 145 1335 155 1355
rect 175 1335 185 1355
rect 145 1325 185 1335
rect -185 1315 -145 1325
rect -185 805 -165 1315
rect -125 1090 -60 1100
rect -125 1070 -115 1090
rect -70 1070 -60 1090
rect -125 1060 -60 1070
rect 60 1090 125 1100
rect 60 1070 70 1090
rect 115 1070 125 1090
rect 60 1060 125 1070
rect 165 815 185 1325
rect 145 805 185 815
rect -185 795 -145 805
rect -185 775 -175 795
rect -155 775 -145 795
rect 145 785 155 805
rect 175 785 185 805
rect 145 775 185 785
rect 355 1915 375 2290
rect 705 2415 725 2425
rect 895 2455 935 2465
rect 895 2435 905 2455
rect 925 2435 935 2455
rect 895 2425 935 2435
rect 1225 2455 1265 2465
rect 1225 2435 1235 2455
rect 1255 2435 1265 2455
rect 1225 2425 1265 2435
rect 705 2405 800 2415
rect 705 2375 735 2405
rect 790 2375 800 2405
rect 705 2365 800 2375
rect 415 2190 480 2200
rect 415 2170 425 2190
rect 470 2170 480 2190
rect 415 2160 480 2170
rect 600 2190 665 2200
rect 600 2170 610 2190
rect 655 2170 665 2190
rect 600 2160 665 2170
rect 705 1915 725 2365
rect 895 2340 915 2425
rect 820 2330 915 2340
rect 820 2300 830 2330
rect 885 2300 915 2330
rect 820 2290 915 2300
rect 355 1905 395 1915
rect 355 1885 365 1905
rect 385 1885 395 1905
rect 355 1875 395 1885
rect 685 1905 725 1915
rect 685 1885 695 1905
rect 715 1885 725 1905
rect 685 1875 725 1885
rect 355 1365 375 1875
rect 520 1860 560 1870
rect 520 1790 530 1860
rect 550 1790 560 1860
rect 520 1780 560 1790
rect 415 1640 480 1650
rect 415 1620 425 1640
rect 470 1620 480 1640
rect 415 1610 480 1620
rect 600 1640 665 1650
rect 600 1620 610 1640
rect 655 1620 665 1640
rect 600 1610 665 1620
rect 705 1365 725 1875
rect 355 1355 395 1365
rect 355 1335 365 1355
rect 385 1335 395 1355
rect 355 1325 395 1335
rect 685 1355 725 1365
rect 685 1335 695 1355
rect 715 1335 725 1355
rect 685 1325 725 1335
rect 355 815 375 1325
rect 415 1090 480 1100
rect 415 1070 425 1090
rect 470 1070 480 1090
rect 415 1060 480 1070
rect 600 1090 665 1100
rect 600 1070 610 1090
rect 655 1070 665 1090
rect 600 1060 665 1070
rect 705 815 725 1325
rect 355 805 395 815
rect 355 785 365 805
rect 385 785 395 805
rect 355 775 395 785
rect 685 805 725 815
rect 685 785 695 805
rect 715 785 725 805
rect 685 775 725 785
rect 895 1915 915 2290
rect 1245 2415 1265 2425
rect 1435 2455 1475 2465
rect 1435 2435 1445 2455
rect 1465 2435 1475 2455
rect 1435 2425 1475 2435
rect 1765 2455 1805 2465
rect 1765 2435 1775 2455
rect 1795 2435 1805 2455
rect 1765 2425 1805 2435
rect 1245 2405 1340 2415
rect 1245 2375 1275 2405
rect 1330 2375 1340 2405
rect 1245 2365 1340 2375
rect 955 2190 1020 2200
rect 955 2170 965 2190
rect 1010 2170 1020 2190
rect 955 2160 1020 2170
rect 1140 2190 1205 2200
rect 1140 2170 1150 2190
rect 1195 2170 1205 2190
rect 1140 2160 1205 2170
rect 1245 1915 1265 2365
rect 1435 2340 1455 2425
rect 1360 2330 1455 2340
rect 1360 2300 1370 2330
rect 1425 2300 1455 2330
rect 1360 2290 1455 2300
rect 895 1905 935 1915
rect 895 1885 905 1905
rect 925 1885 935 1905
rect 895 1875 935 1885
rect 1225 1905 1265 1915
rect 1225 1885 1235 1905
rect 1255 1885 1265 1905
rect 1225 1875 1265 1885
rect 895 1365 915 1875
rect 1060 1860 1100 1870
rect 1060 1790 1070 1860
rect 1090 1790 1100 1860
rect 1060 1780 1100 1790
rect 955 1640 1020 1650
rect 955 1620 965 1640
rect 1010 1620 1020 1640
rect 955 1610 1020 1620
rect 1140 1640 1205 1650
rect 1140 1620 1150 1640
rect 1195 1620 1205 1640
rect 1140 1610 1205 1620
rect 1245 1365 1265 1875
rect 895 1355 935 1365
rect 895 1335 905 1355
rect 925 1335 935 1355
rect 895 1325 935 1335
rect 1225 1355 1265 1365
rect 1225 1335 1235 1355
rect 1255 1335 1265 1355
rect 1225 1325 1265 1335
rect 895 815 915 1325
rect 955 1090 1020 1100
rect 955 1070 965 1090
rect 1010 1070 1020 1090
rect 955 1060 1020 1070
rect 1140 1090 1205 1100
rect 1140 1070 1150 1090
rect 1195 1070 1205 1090
rect 1140 1060 1205 1070
rect 1245 815 1265 1325
rect 895 805 935 815
rect 895 785 905 805
rect 925 785 935 805
rect 895 775 935 785
rect 1225 805 1265 815
rect 1225 785 1235 805
rect 1255 785 1265 805
rect 1225 775 1265 785
rect 1435 1915 1455 2290
rect 1785 2415 1805 2425
rect 1975 2455 2015 2465
rect 1975 2435 1985 2455
rect 2005 2435 2015 2455
rect 1975 2425 2015 2435
rect 2305 2455 2345 2465
rect 2305 2435 2315 2455
rect 2335 2435 2345 2455
rect 2305 2425 2345 2435
rect 1785 2405 1880 2415
rect 1785 2375 1815 2405
rect 1870 2375 1880 2405
rect 1785 2365 1880 2375
rect 1495 2190 1560 2200
rect 1495 2170 1505 2190
rect 1550 2170 1560 2190
rect 1495 2160 1560 2170
rect 1680 2190 1745 2200
rect 1680 2170 1690 2190
rect 1735 2170 1745 2190
rect 1680 2160 1745 2170
rect 1785 1915 1805 2365
rect 1975 2340 1995 2425
rect 1900 2330 1995 2340
rect 1900 2300 1910 2330
rect 1965 2300 1995 2330
rect 1900 2290 1995 2300
rect 1435 1905 1475 1915
rect 1435 1885 1445 1905
rect 1465 1885 1475 1905
rect 1435 1875 1475 1885
rect 1765 1905 1805 1915
rect 1765 1885 1775 1905
rect 1795 1885 1805 1905
rect 1765 1875 1805 1885
rect 1435 1365 1455 1875
rect 1600 1860 1640 1870
rect 1600 1790 1610 1860
rect 1630 1790 1640 1860
rect 1600 1780 1640 1790
rect 1495 1640 1560 1650
rect 1495 1620 1505 1640
rect 1550 1620 1560 1640
rect 1495 1610 1560 1620
rect 1680 1640 1745 1650
rect 1680 1620 1690 1640
rect 1735 1620 1745 1640
rect 1680 1610 1745 1620
rect 1785 1365 1805 1875
rect 1435 1355 1475 1365
rect 1435 1335 1445 1355
rect 1465 1335 1475 1355
rect 1435 1325 1475 1335
rect 1765 1355 1805 1365
rect 1765 1335 1775 1355
rect 1795 1335 1805 1355
rect 1765 1325 1805 1335
rect 1435 815 1455 1325
rect 1495 1090 1560 1100
rect 1495 1070 1505 1090
rect 1550 1070 1560 1090
rect 1495 1060 1560 1070
rect 1680 1090 1745 1100
rect 1680 1070 1690 1090
rect 1735 1070 1745 1090
rect 1680 1060 1745 1070
rect 1785 815 1805 1325
rect 1435 805 1475 815
rect 1435 785 1445 805
rect 1465 785 1475 805
rect 1435 775 1475 785
rect 1765 805 1805 815
rect 1765 785 1775 805
rect 1795 785 1805 805
rect 1765 775 1805 785
rect 1975 1915 1995 2290
rect 2325 2415 2345 2425
rect 2515 2455 2555 2465
rect 2515 2435 2525 2455
rect 2545 2435 2555 2455
rect 2515 2425 2555 2435
rect 2845 2455 2885 2465
rect 2845 2435 2855 2455
rect 2875 2435 2885 2455
rect 2845 2425 2885 2435
rect 2325 2405 2420 2415
rect 2325 2375 2355 2405
rect 2410 2375 2420 2405
rect 2325 2365 2420 2375
rect 2035 2190 2100 2200
rect 2035 2170 2045 2190
rect 2090 2170 2100 2190
rect 2035 2160 2100 2170
rect 2220 2190 2285 2200
rect 2220 2170 2230 2190
rect 2275 2170 2285 2190
rect 2220 2160 2285 2170
rect 2325 1915 2345 2365
rect 2515 2340 2535 2425
rect 2440 2330 2535 2340
rect 2440 2300 2450 2330
rect 2505 2300 2535 2330
rect 2440 2290 2535 2300
rect 1975 1905 2015 1915
rect 1975 1885 1985 1905
rect 2005 1885 2015 1905
rect 1975 1875 2015 1885
rect 2305 1905 2345 1915
rect 2305 1885 2315 1905
rect 2335 1885 2345 1905
rect 2305 1875 2345 1885
rect 1975 1365 1995 1875
rect 2140 1860 2180 1870
rect 2140 1790 2150 1860
rect 2170 1790 2180 1860
rect 2140 1780 2180 1790
rect 2035 1640 2100 1650
rect 2035 1620 2045 1640
rect 2090 1620 2100 1640
rect 2035 1610 2100 1620
rect 2220 1640 2285 1650
rect 2220 1620 2230 1640
rect 2275 1620 2285 1640
rect 2220 1610 2285 1620
rect 2325 1365 2345 1875
rect 1975 1355 2015 1365
rect 1975 1335 1985 1355
rect 2005 1335 2015 1355
rect 1975 1325 2015 1335
rect 2305 1355 2345 1365
rect 2305 1335 2315 1355
rect 2335 1335 2345 1355
rect 2305 1325 2345 1335
rect 1975 815 1995 1325
rect 2035 1090 2100 1100
rect 2035 1070 2045 1090
rect 2090 1070 2100 1090
rect 2035 1060 2100 1070
rect 2220 1090 2285 1100
rect 2220 1070 2230 1090
rect 2275 1070 2285 1090
rect 2220 1060 2285 1070
rect 2325 815 2345 1325
rect 1975 805 2015 815
rect 1975 785 1985 805
rect 2005 785 2015 805
rect 1975 775 2015 785
rect 2305 805 2345 815
rect 2305 785 2315 805
rect 2335 785 2345 805
rect 2305 775 2345 785
rect 2515 1915 2535 2290
rect 2865 2415 2885 2425
rect 3055 2455 3095 2465
rect 3055 2435 3065 2455
rect 3085 2435 3095 2455
rect 3055 2425 3095 2435
rect 3385 2455 3425 2465
rect 3385 2435 3395 2455
rect 3415 2435 3425 2455
rect 3385 2425 3425 2435
rect 2865 2405 2960 2415
rect 2865 2375 2895 2405
rect 2950 2375 2960 2405
rect 2865 2365 2960 2375
rect 2575 2190 2640 2200
rect 2575 2170 2585 2190
rect 2630 2170 2640 2190
rect 2575 2160 2640 2170
rect 2760 2190 2825 2200
rect 2760 2170 2770 2190
rect 2815 2170 2825 2190
rect 2760 2160 2825 2170
rect 2865 1915 2885 2365
rect 3055 2340 3075 2425
rect 2980 2330 3075 2340
rect 2980 2300 2990 2330
rect 3045 2300 3075 2330
rect 2980 2290 3075 2300
rect 2515 1905 2555 1915
rect 2515 1885 2525 1905
rect 2545 1885 2555 1905
rect 2515 1875 2555 1885
rect 2845 1905 2885 1915
rect 2845 1885 2855 1905
rect 2875 1885 2885 1905
rect 2845 1875 2885 1885
rect 2515 1365 2535 1875
rect 2680 1860 2720 1870
rect 2680 1790 2690 1860
rect 2710 1790 2720 1860
rect 2680 1780 2720 1790
rect 2575 1640 2640 1650
rect 2575 1620 2585 1640
rect 2630 1620 2640 1640
rect 2575 1610 2640 1620
rect 2760 1640 2825 1650
rect 2760 1620 2770 1640
rect 2815 1620 2825 1640
rect 2760 1610 2825 1620
rect 2865 1365 2885 1875
rect 2515 1355 2555 1365
rect 2515 1335 2525 1355
rect 2545 1335 2555 1355
rect 2515 1325 2555 1335
rect 2845 1355 2885 1365
rect 2845 1335 2855 1355
rect 2875 1335 2885 1355
rect 2845 1325 2885 1335
rect 2515 815 2535 1325
rect 2575 1090 2640 1100
rect 2575 1070 2585 1090
rect 2630 1070 2640 1090
rect 2575 1060 2640 1070
rect 2760 1090 2825 1100
rect 2760 1070 2770 1090
rect 2815 1070 2825 1090
rect 2760 1060 2825 1070
rect 2865 815 2885 1325
rect 2515 805 2555 815
rect 2515 785 2525 805
rect 2545 785 2555 805
rect 2515 775 2555 785
rect 2845 805 2885 815
rect 2845 785 2855 805
rect 2875 785 2885 805
rect 2845 775 2885 785
rect 3055 1915 3075 2290
rect 3115 2190 3180 2200
rect 3115 2170 3125 2190
rect 3170 2170 3180 2190
rect 3115 2160 3180 2170
rect 3300 2190 3365 2200
rect 3300 2170 3310 2190
rect 3355 2170 3365 2190
rect 3300 2160 3365 2170
rect 3405 1915 3425 2425
rect 3055 1905 3095 1915
rect 3055 1885 3065 1905
rect 3085 1885 3095 1905
rect 3055 1875 3095 1885
rect 3385 1905 3425 1915
rect 3385 1885 3395 1905
rect 3415 1885 3425 1905
rect 3385 1875 3425 1885
rect 3055 1365 3075 1875
rect 3220 1860 3260 1870
rect 3220 1790 3230 1860
rect 3250 1790 3260 1860
rect 3220 1780 3260 1790
rect 3115 1640 3180 1650
rect 3115 1620 3125 1640
rect 3170 1620 3180 1640
rect 3115 1610 3180 1620
rect 3300 1640 3365 1650
rect 3300 1620 3310 1640
rect 3355 1620 3365 1640
rect 3300 1610 3365 1620
rect 3405 1365 3425 1875
rect 3055 1355 3095 1365
rect 3055 1335 3065 1355
rect 3085 1335 3095 1355
rect 3055 1325 3095 1335
rect 3385 1355 3425 1365
rect 3385 1335 3395 1355
rect 3415 1335 3425 1355
rect 3385 1325 3425 1335
rect 3055 815 3075 1325
rect 3115 1090 3180 1100
rect 3115 1070 3125 1090
rect 3170 1070 3180 1090
rect 3115 1060 3180 1070
rect 3300 1090 3365 1100
rect 3300 1070 3310 1090
rect 3355 1070 3365 1090
rect 3300 1060 3365 1070
rect 3405 815 3425 1325
rect 3055 805 3095 815
rect 3055 785 3065 805
rect 3085 785 3095 805
rect 3055 775 3095 785
rect 3385 805 3425 815
rect 3385 785 3395 805
rect 3415 785 3425 805
rect 3385 775 3425 785
rect -185 765 -145 775
rect -125 540 -60 550
rect -125 520 -115 540
rect -70 520 -60 540
rect -125 510 -60 520
rect 60 540 125 550
rect 60 520 70 540
rect 115 520 125 540
rect 60 510 125 520
rect 415 540 480 550
rect 415 520 425 540
rect 470 520 480 540
rect 415 510 480 520
rect 600 540 665 550
rect 600 520 610 540
rect 655 520 665 540
rect 600 510 665 520
rect 955 540 1020 550
rect 955 520 965 540
rect 1010 520 1020 540
rect 955 510 1020 520
rect 1140 540 1205 550
rect 1140 520 1150 540
rect 1195 520 1205 540
rect 1140 510 1205 520
rect 1495 540 1560 550
rect 1495 520 1505 540
rect 1550 520 1560 540
rect 1495 510 1560 520
rect 1680 540 1745 550
rect 1680 520 1690 540
rect 1735 520 1745 540
rect 1680 510 1745 520
rect 2035 540 2100 550
rect 2035 520 2045 540
rect 2090 520 2100 540
rect 2035 510 2100 520
rect 2220 540 2285 550
rect 2220 520 2230 540
rect 2275 520 2285 540
rect 2220 510 2285 520
rect 2575 540 2640 550
rect 2575 520 2585 540
rect 2630 520 2640 540
rect 2575 510 2640 520
rect 2760 540 2825 550
rect 2760 520 2770 540
rect 2815 520 2825 540
rect 2760 510 2825 520
rect 3115 540 3180 550
rect 3115 520 3125 540
rect 3170 520 3180 540
rect 3115 510 3180 520
rect 3300 540 3365 550
rect 3300 520 3310 540
rect 3355 520 3365 540
rect 3300 510 3365 520
rect -125 505 -105 510
rect 415 505 435 510
rect 955 505 975 510
rect 1495 505 1515 510
rect 2035 505 2055 510
rect 2575 505 2595 510
rect 3115 505 3135 510
rect -125 420 -105 425
rect 60 420 80 425
rect 415 420 435 425
rect 600 420 620 425
rect 955 420 975 425
rect 1140 420 1160 425
rect 1495 420 1515 425
rect 1680 420 1700 425
rect 2035 420 2055 425
rect 2220 420 2240 425
rect 2575 420 2595 425
rect 2760 420 2780 425
rect 3115 420 3135 425
rect 3300 420 3320 425
rect -125 410 -60 420
rect -125 390 -115 410
rect -70 390 -60 410
rect -125 380 -60 390
rect 60 410 250 420
rect 60 390 70 410
rect 115 400 250 410
rect 115 390 125 400
rect 60 380 125 390
rect -185 120 -145 130
rect -185 100 -175 120
rect -155 100 -145 120
rect -185 90 -145 100
rect 145 120 185 130
rect 145 100 155 120
rect 175 100 185 120
rect 145 90 185 100
rect -185 -420 -165 90
rect -125 -140 -60 -130
rect -125 -160 -115 -140
rect -70 -160 -60 -140
rect -125 -170 -60 -160
rect 60 -140 125 -130
rect 60 -160 70 -140
rect 115 -160 125 -140
rect 60 -170 125 -160
rect 165 -420 185 90
rect -185 -430 -145 -420
rect -185 -450 -175 -430
rect -155 -450 -145 -430
rect -185 -460 -145 -450
rect 145 -430 185 -420
rect 145 -450 155 -430
rect 175 -450 185 -430
rect 145 -460 185 -450
rect -185 -970 -165 -460
rect -125 -690 -60 -680
rect -125 -710 -115 -690
rect -70 -710 -60 -690
rect -125 -720 -60 -710
rect 60 -690 125 -680
rect 60 -710 70 -690
rect 115 -710 125 -690
rect 60 -720 125 -710
rect 165 -970 185 -460
rect -185 -980 -145 -970
rect -185 -1000 -175 -980
rect -155 -1000 -145 -980
rect -185 -1010 -145 -1000
rect 145 -980 185 -970
rect 145 -1000 155 -980
rect 175 -1000 185 -980
rect 145 -1010 185 -1000
rect -185 -1520 -165 -1010
rect -20 -1020 20 -1010
rect -20 -1090 -10 -1020
rect 10 -1090 20 -1020
rect -20 -1100 20 -1090
rect -125 -1240 -60 -1230
rect -125 -1260 -115 -1240
rect -70 -1260 -60 -1240
rect -125 -1270 -60 -1260
rect 60 -1240 125 -1230
rect 60 -1260 70 -1240
rect 115 -1260 125 -1240
rect 60 -1270 125 -1260
rect 165 -1520 185 -1010
rect -185 -1530 -145 -1520
rect -185 -1550 -175 -1530
rect -155 -1550 -145 -1530
rect -185 -1560 -145 -1550
rect 145 -1530 185 -1520
rect 145 -1550 155 -1530
rect 175 -1550 185 -1530
rect 145 -1560 185 -1550
rect 230 -1780 250 400
rect 415 410 480 420
rect 415 390 425 410
rect 470 390 480 410
rect 415 380 480 390
rect 600 410 795 420
rect 600 390 610 410
rect 655 400 795 410
rect 655 390 665 400
rect 600 380 665 390
rect 355 120 395 130
rect 355 100 365 120
rect 385 100 395 120
rect 355 90 395 100
rect 685 120 725 130
rect 685 100 695 120
rect 715 100 725 120
rect 685 90 725 100
rect 355 -420 375 90
rect 415 -140 480 -130
rect 415 -160 425 -140
rect 470 -160 480 -140
rect 415 -170 480 -160
rect 600 -140 665 -130
rect 600 -160 610 -140
rect 655 -160 665 -140
rect 600 -170 665 -160
rect 705 -420 725 90
rect 355 -430 395 -420
rect 355 -450 365 -430
rect 385 -450 395 -430
rect 355 -460 395 -450
rect 685 -430 725 -420
rect 685 -450 695 -430
rect 715 -450 725 -430
rect 685 -460 725 -450
rect 355 -970 375 -460
rect 415 -690 480 -680
rect 415 -710 425 -690
rect 470 -710 480 -690
rect 415 -720 480 -710
rect 600 -690 665 -680
rect 600 -710 610 -690
rect 655 -710 665 -690
rect 600 -720 665 -710
rect 705 -970 725 -460
rect 355 -980 395 -970
rect 355 -1000 365 -980
rect 385 -1000 395 -980
rect 355 -1010 395 -1000
rect 685 -980 725 -970
rect 685 -1000 695 -980
rect 715 -1000 725 -980
rect 685 -1010 725 -1000
rect 355 -1520 375 -1010
rect 520 -1020 560 -1010
rect 520 -1090 530 -1020
rect 550 -1090 560 -1020
rect 520 -1100 560 -1090
rect 415 -1240 480 -1230
rect 415 -1260 425 -1240
rect 470 -1260 480 -1240
rect 415 -1270 480 -1260
rect 600 -1240 665 -1230
rect 600 -1260 610 -1240
rect 655 -1260 665 -1240
rect 600 -1270 665 -1260
rect 705 -1520 725 -1010
rect 355 -1530 395 -1520
rect 355 -1550 365 -1530
rect 385 -1550 395 -1530
rect 355 -1560 395 -1550
rect 685 -1530 725 -1520
rect 685 -1550 695 -1530
rect 715 -1550 725 -1530
rect 685 -1560 725 -1550
rect 775 -1780 795 400
rect 955 410 1020 420
rect 955 390 965 410
rect 1010 390 1020 410
rect 955 380 1020 390
rect 1140 410 1335 420
rect 1140 390 1150 410
rect 1195 400 1335 410
rect 1195 390 1205 400
rect 1140 380 1205 390
rect 895 120 935 130
rect 895 100 905 120
rect 925 100 935 120
rect 895 90 935 100
rect 1225 120 1265 130
rect 1225 100 1235 120
rect 1255 100 1265 120
rect 1225 90 1265 100
rect 895 -420 915 90
rect 955 -140 1020 -130
rect 955 -160 965 -140
rect 1010 -160 1020 -140
rect 955 -170 1020 -160
rect 1140 -140 1205 -130
rect 1140 -160 1150 -140
rect 1195 -160 1205 -140
rect 1140 -170 1205 -160
rect 1245 -420 1265 90
rect 895 -430 935 -420
rect 895 -450 905 -430
rect 925 -450 935 -430
rect 895 -460 935 -450
rect 1225 -430 1265 -420
rect 1225 -450 1235 -430
rect 1255 -450 1265 -430
rect 1225 -460 1265 -450
rect 895 -970 915 -460
rect 955 -690 1020 -680
rect 955 -710 965 -690
rect 1010 -710 1020 -690
rect 955 -720 1020 -710
rect 1140 -690 1205 -680
rect 1140 -710 1150 -690
rect 1195 -710 1205 -690
rect 1140 -720 1205 -710
rect 1245 -970 1265 -460
rect 895 -980 935 -970
rect 895 -1000 905 -980
rect 925 -1000 935 -980
rect 895 -1010 935 -1000
rect 1225 -980 1265 -970
rect 1225 -1000 1235 -980
rect 1255 -1000 1265 -980
rect 1225 -1010 1265 -1000
rect 895 -1520 915 -1010
rect 1060 -1020 1100 -1010
rect 1060 -1090 1070 -1020
rect 1090 -1090 1100 -1020
rect 1060 -1100 1100 -1090
rect 955 -1240 1020 -1230
rect 955 -1260 965 -1240
rect 1010 -1260 1020 -1240
rect 955 -1270 1020 -1260
rect 1140 -1240 1205 -1230
rect 1140 -1260 1150 -1240
rect 1195 -1260 1205 -1240
rect 1140 -1270 1205 -1260
rect 1245 -1520 1265 -1010
rect 895 -1530 935 -1520
rect 895 -1550 905 -1530
rect 925 -1550 935 -1530
rect 895 -1560 935 -1550
rect 1225 -1530 1265 -1520
rect 1225 -1550 1235 -1530
rect 1255 -1550 1265 -1530
rect 1225 -1560 1265 -1550
rect 1315 -1780 1335 400
rect 1495 410 1560 420
rect 1495 390 1505 410
rect 1550 390 1560 410
rect 1495 380 1560 390
rect 1680 410 1875 420
rect 1680 390 1690 410
rect 1735 400 1875 410
rect 1735 390 1745 400
rect 1680 380 1745 390
rect 1435 120 1475 130
rect 1435 100 1445 120
rect 1465 100 1475 120
rect 1435 90 1475 100
rect 1765 120 1805 130
rect 1765 100 1775 120
rect 1795 100 1805 120
rect 1765 90 1805 100
rect 1435 -420 1455 90
rect 1495 -140 1560 -130
rect 1495 -160 1505 -140
rect 1550 -160 1560 -140
rect 1495 -170 1560 -160
rect 1680 -140 1745 -130
rect 1680 -160 1690 -140
rect 1735 -160 1745 -140
rect 1680 -170 1745 -160
rect 1785 -420 1805 90
rect 1435 -430 1475 -420
rect 1435 -450 1445 -430
rect 1465 -450 1475 -430
rect 1435 -460 1475 -450
rect 1765 -430 1805 -420
rect 1765 -450 1775 -430
rect 1795 -450 1805 -430
rect 1765 -460 1805 -450
rect 1435 -970 1455 -460
rect 1495 -690 1560 -680
rect 1495 -710 1505 -690
rect 1550 -710 1560 -690
rect 1495 -720 1560 -710
rect 1680 -690 1745 -680
rect 1680 -710 1690 -690
rect 1735 -710 1745 -690
rect 1680 -720 1745 -710
rect 1785 -970 1805 -460
rect 1435 -980 1475 -970
rect 1435 -1000 1445 -980
rect 1465 -1000 1475 -980
rect 1435 -1010 1475 -1000
rect 1765 -980 1805 -970
rect 1765 -1000 1775 -980
rect 1795 -1000 1805 -980
rect 1765 -1010 1805 -1000
rect 1435 -1520 1455 -1010
rect 1600 -1020 1640 -1010
rect 1600 -1090 1610 -1020
rect 1630 -1090 1640 -1020
rect 1600 -1100 1640 -1090
rect 1495 -1240 1560 -1230
rect 1495 -1260 1505 -1240
rect 1550 -1260 1560 -1240
rect 1495 -1270 1560 -1260
rect 1680 -1240 1745 -1230
rect 1680 -1260 1690 -1240
rect 1735 -1260 1745 -1240
rect 1680 -1270 1745 -1260
rect 1785 -1520 1805 -1010
rect 1435 -1530 1475 -1520
rect 1435 -1550 1445 -1530
rect 1465 -1550 1475 -1530
rect 1435 -1560 1475 -1550
rect 1765 -1530 1805 -1520
rect 1765 -1550 1775 -1530
rect 1795 -1550 1805 -1530
rect 1765 -1560 1805 -1550
rect 1855 -1780 1875 400
rect 2035 410 2100 420
rect 2035 390 2045 410
rect 2090 390 2100 410
rect 2035 380 2100 390
rect 2220 410 2415 420
rect 2220 390 2230 410
rect 2275 400 2415 410
rect 2275 390 2285 400
rect 2220 380 2285 390
rect 1975 120 2015 130
rect 1975 100 1985 120
rect 2005 100 2015 120
rect 1975 90 2015 100
rect 2305 120 2345 130
rect 2305 100 2315 120
rect 2335 100 2345 120
rect 2305 90 2345 100
rect 1975 -420 1995 90
rect 2035 -140 2100 -130
rect 2035 -160 2045 -140
rect 2090 -160 2100 -140
rect 2035 -170 2100 -160
rect 2220 -140 2285 -130
rect 2220 -160 2230 -140
rect 2275 -160 2285 -140
rect 2220 -170 2285 -160
rect 2325 -420 2345 90
rect 1975 -430 2015 -420
rect 1975 -450 1985 -430
rect 2005 -450 2015 -430
rect 1975 -460 2015 -450
rect 2305 -430 2345 -420
rect 2305 -450 2315 -430
rect 2335 -450 2345 -430
rect 2305 -460 2345 -450
rect 1975 -970 1995 -460
rect 2035 -690 2100 -680
rect 2035 -710 2045 -690
rect 2090 -710 2100 -690
rect 2035 -720 2100 -710
rect 2220 -690 2285 -680
rect 2220 -710 2230 -690
rect 2275 -710 2285 -690
rect 2220 -720 2285 -710
rect 2325 -970 2345 -460
rect 1975 -980 2015 -970
rect 1975 -1000 1985 -980
rect 2005 -1000 2015 -980
rect 1975 -1010 2015 -1000
rect 2305 -980 2345 -970
rect 2305 -1000 2315 -980
rect 2335 -1000 2345 -980
rect 2305 -1010 2345 -1000
rect 1975 -1520 1995 -1010
rect 2140 -1020 2180 -1010
rect 2140 -1090 2150 -1020
rect 2170 -1090 2180 -1020
rect 2140 -1100 2180 -1090
rect 2035 -1240 2100 -1230
rect 2035 -1260 2045 -1240
rect 2090 -1260 2100 -1240
rect 2035 -1270 2100 -1260
rect 2220 -1240 2285 -1230
rect 2220 -1260 2230 -1240
rect 2275 -1260 2285 -1240
rect 2220 -1270 2285 -1260
rect 2325 -1520 2345 -1010
rect 1975 -1530 2015 -1520
rect 1975 -1550 1985 -1530
rect 2005 -1550 2015 -1530
rect 1975 -1560 2015 -1550
rect 2305 -1530 2345 -1520
rect 2305 -1550 2315 -1530
rect 2335 -1550 2345 -1530
rect 2305 -1560 2345 -1550
rect 2395 -1780 2415 400
rect 2575 410 2640 420
rect 2575 390 2585 410
rect 2630 390 2640 410
rect 2575 380 2640 390
rect 2760 410 2955 420
rect 2760 390 2770 410
rect 2815 400 2955 410
rect 2815 390 2825 400
rect 2760 380 2825 390
rect 2515 120 2555 130
rect 2515 100 2525 120
rect 2545 100 2555 120
rect 2515 90 2555 100
rect 2845 120 2885 130
rect 2845 100 2855 120
rect 2875 100 2885 120
rect 2845 90 2885 100
rect 2515 -420 2535 90
rect 2575 -140 2640 -130
rect 2575 -160 2585 -140
rect 2630 -160 2640 -140
rect 2575 -170 2640 -160
rect 2760 -140 2825 -130
rect 2760 -160 2770 -140
rect 2815 -160 2825 -140
rect 2760 -170 2825 -160
rect 2865 -420 2885 90
rect 2515 -430 2555 -420
rect 2515 -450 2525 -430
rect 2545 -450 2555 -430
rect 2515 -460 2555 -450
rect 2845 -430 2885 -420
rect 2845 -450 2855 -430
rect 2875 -450 2885 -430
rect 2845 -460 2885 -450
rect 2515 -970 2535 -460
rect 2575 -690 2640 -680
rect 2575 -710 2585 -690
rect 2630 -710 2640 -690
rect 2575 -720 2640 -710
rect 2760 -690 2825 -680
rect 2760 -710 2770 -690
rect 2815 -710 2825 -690
rect 2760 -720 2825 -710
rect 2865 -970 2885 -460
rect 2515 -980 2555 -970
rect 2515 -1000 2525 -980
rect 2545 -1000 2555 -980
rect 2515 -1010 2555 -1000
rect 2845 -980 2885 -970
rect 2845 -1000 2855 -980
rect 2875 -1000 2885 -980
rect 2845 -1010 2885 -1000
rect 2515 -1520 2535 -1010
rect 2680 -1020 2720 -1010
rect 2680 -1090 2690 -1020
rect 2710 -1090 2720 -1020
rect 2680 -1100 2720 -1090
rect 2575 -1240 2640 -1230
rect 2575 -1260 2585 -1240
rect 2630 -1260 2640 -1240
rect 2575 -1270 2640 -1260
rect 2760 -1240 2825 -1230
rect 2760 -1260 2770 -1240
rect 2815 -1260 2825 -1240
rect 2760 -1270 2825 -1260
rect 2865 -1520 2885 -1010
rect 2515 -1530 2555 -1520
rect 2515 -1550 2525 -1530
rect 2545 -1550 2555 -1530
rect 2515 -1560 2555 -1550
rect 2845 -1530 2885 -1520
rect 2845 -1550 2855 -1530
rect 2875 -1550 2885 -1530
rect 2845 -1560 2885 -1550
rect 2935 -1780 2955 400
rect 3115 410 3180 420
rect 3115 390 3125 410
rect 3170 390 3180 410
rect 3115 380 3180 390
rect 3300 410 3530 420
rect 3300 390 3310 410
rect 3355 400 3530 410
rect 3355 390 3365 400
rect 3300 380 3365 390
rect 3055 120 3095 130
rect 3055 100 3065 120
rect 3085 100 3095 120
rect 3055 90 3095 100
rect 3385 120 3425 130
rect 3385 100 3395 120
rect 3415 100 3425 120
rect 3385 90 3425 100
rect 3055 -420 3075 90
rect 3115 -140 3180 -130
rect 3115 -160 3125 -140
rect 3170 -160 3180 -140
rect 3115 -170 3180 -160
rect 3300 -140 3365 -130
rect 3300 -160 3310 -140
rect 3355 -160 3365 -140
rect 3300 -170 3365 -160
rect 3405 -420 3425 90
rect 3055 -430 3095 -420
rect 3055 -450 3065 -430
rect 3085 -450 3095 -430
rect 3055 -460 3095 -450
rect 3385 -430 3425 -420
rect 3385 -450 3395 -430
rect 3415 -450 3425 -430
rect 3385 -460 3425 -450
rect 3055 -970 3075 -460
rect 3115 -690 3180 -680
rect 3115 -710 3125 -690
rect 3170 -710 3180 -690
rect 3115 -720 3180 -710
rect 3300 -690 3365 -680
rect 3300 -710 3310 -690
rect 3355 -710 3365 -690
rect 3300 -720 3365 -710
rect 3405 -970 3425 -460
rect 3055 -980 3095 -970
rect 3055 -1000 3065 -980
rect 3085 -1000 3095 -980
rect 3055 -1010 3095 -1000
rect 3385 -980 3425 -970
rect 3385 -1000 3395 -980
rect 3415 -1000 3425 -980
rect 3385 -1010 3425 -1000
rect 3055 -1520 3075 -1010
rect 3220 -1020 3260 -1010
rect 3220 -1090 3230 -1020
rect 3250 -1090 3260 -1020
rect 3220 -1100 3260 -1090
rect 3115 -1240 3180 -1230
rect 3115 -1260 3125 -1240
rect 3170 -1260 3180 -1240
rect 3115 -1270 3180 -1260
rect 3300 -1240 3365 -1230
rect 3300 -1260 3310 -1240
rect 3355 -1260 3365 -1240
rect 3300 -1270 3365 -1260
rect 3405 -1520 3425 -1010
rect 3055 -1530 3095 -1520
rect 3055 -1550 3065 -1530
rect 3085 -1550 3095 -1530
rect 3055 -1560 3095 -1550
rect 3385 -1530 3425 -1520
rect 3385 -1550 3395 -1530
rect 3415 -1550 3425 -1530
rect 3385 -1560 3425 -1550
rect 3510 -1780 3530 400
rect 3655 410 3720 420
rect 3655 390 3665 410
rect 3710 390 3720 410
rect 3655 380 3720 390
rect 3740 120 3780 130
rect 3740 100 3750 120
rect 3770 100 3780 120
rect 3740 90 3780 100
rect 3655 -140 3720 -130
rect 3655 -160 3665 -140
rect 3710 -160 3720 -140
rect 3655 -170 3720 -160
rect 3760 -420 3780 90
rect 3740 -430 3780 -420
rect 3740 -450 3750 -430
rect 3770 -450 3780 -430
rect 3740 -460 3780 -450
rect 3655 -690 3720 -680
rect 3655 -710 3665 -690
rect 3710 -710 3720 -690
rect 3655 -720 3720 -710
rect 3760 -970 3780 -460
rect 3740 -980 3780 -970
rect 3740 -1000 3750 -980
rect 3770 -1000 3780 -980
rect 3740 -1010 3780 -1000
rect 3655 -1240 3720 -1230
rect 3655 -1260 3665 -1240
rect 3710 -1260 3720 -1240
rect 3655 -1270 3720 -1260
rect 3760 -1520 3780 -1010
rect 3740 -1530 3780 -1520
rect 3740 -1550 3750 -1530
rect 3770 -1550 3780 -1530
rect 3740 -1560 3780 -1550
rect -125 -1790 -60 -1780
rect -125 -1810 -115 -1790
rect -70 -1810 -60 -1790
rect -125 -1820 -60 -1810
rect 60 -1790 125 -1780
rect 60 -1810 70 -1790
rect 115 -1810 125 -1790
rect 230 -1790 480 -1780
rect 230 -1800 425 -1790
rect 60 -1820 125 -1810
rect 415 -1810 425 -1800
rect 470 -1810 480 -1790
rect 415 -1820 480 -1810
rect 600 -1790 665 -1780
rect 600 -1810 610 -1790
rect 655 -1810 665 -1790
rect 775 -1790 1020 -1780
rect 775 -1800 965 -1790
rect 600 -1820 665 -1810
rect 955 -1810 965 -1800
rect 1010 -1810 1020 -1790
rect 955 -1820 1020 -1810
rect 1140 -1790 1205 -1780
rect 1140 -1810 1150 -1790
rect 1195 -1810 1205 -1790
rect 1315 -1790 1560 -1780
rect 1315 -1800 1505 -1790
rect 1140 -1820 1205 -1810
rect 1495 -1810 1505 -1800
rect 1550 -1810 1560 -1790
rect 1495 -1820 1560 -1810
rect 1680 -1790 1745 -1780
rect 1680 -1810 1690 -1790
rect 1735 -1810 1745 -1790
rect 1855 -1790 2100 -1780
rect 1855 -1800 2045 -1790
rect 1680 -1820 1745 -1810
rect 2035 -1810 2045 -1800
rect 2090 -1810 2100 -1790
rect 2035 -1820 2100 -1810
rect 2220 -1790 2285 -1780
rect 2220 -1810 2230 -1790
rect 2275 -1810 2285 -1790
rect 2395 -1790 2640 -1780
rect 2395 -1800 2585 -1790
rect 2220 -1820 2285 -1810
rect 2575 -1810 2585 -1800
rect 2630 -1810 2640 -1790
rect 2575 -1820 2640 -1810
rect 2760 -1790 2825 -1780
rect 2760 -1810 2770 -1790
rect 2815 -1810 2825 -1790
rect 2935 -1790 3180 -1780
rect 2935 -1800 3125 -1790
rect 2760 -1820 2825 -1810
rect 3115 -1810 3125 -1800
rect 3170 -1810 3180 -1790
rect 3115 -1820 3180 -1810
rect 3300 -1790 3365 -1780
rect 3300 -1810 3310 -1790
rect 3355 -1810 3365 -1790
rect 3510 -1790 3720 -1780
rect 3510 -1800 3665 -1790
rect 3300 -1820 3365 -1810
rect 3655 -1810 3665 -1800
rect 3710 -1810 3720 -1790
rect 3655 -1820 3720 -1810
rect -185 -2060 -145 -2050
rect -185 -2080 -175 -2060
rect -155 -2070 -145 -2060
rect 145 -2060 185 -2050
rect 145 -2070 155 -2060
rect -155 -2080 155 -2070
rect 175 -2070 185 -2060
rect 500 -2060 540 -2050
rect 500 -2070 510 -2060
rect 175 -2080 510 -2070
rect 530 -2070 540 -2060
rect 685 -2060 725 -2050
rect 685 -2070 695 -2060
rect 530 -2080 695 -2070
rect 715 -2070 725 -2060
rect 1040 -2060 1080 -2050
rect 1040 -2070 1050 -2060
rect 715 -2080 1050 -2070
rect 1070 -2070 1080 -2060
rect 1225 -2060 1265 -2050
rect 1225 -2070 1235 -2060
rect 1070 -2080 1235 -2070
rect 1255 -2070 1265 -2060
rect 1580 -2060 1620 -2050
rect 1580 -2070 1590 -2060
rect 1255 -2080 1590 -2070
rect 1610 -2070 1620 -2060
rect 1765 -2060 1805 -2050
rect 1765 -2070 1775 -2060
rect 1610 -2080 1775 -2070
rect 1795 -2070 1805 -2060
rect 2120 -2060 2160 -2050
rect 2120 -2070 2130 -2060
rect 1795 -2080 2130 -2070
rect 2150 -2070 2160 -2060
rect 2305 -2060 2345 -2050
rect 2305 -2070 2315 -2060
rect 2150 -2080 2315 -2070
rect 2335 -2070 2345 -2060
rect 2660 -2060 2700 -2050
rect 2660 -2070 2670 -2060
rect 2335 -2080 2670 -2070
rect 2690 -2070 2700 -2060
rect 2845 -2060 2885 -2050
rect 2845 -2070 2855 -2060
rect 2690 -2080 2855 -2070
rect 2875 -2070 2885 -2060
rect 3200 -2060 3240 -2050
rect 3200 -2070 3210 -2060
rect 2875 -2080 3210 -2070
rect 3230 -2070 3240 -2060
rect 3385 -2060 3425 -2050
rect 3385 -2070 3395 -2060
rect 3230 -2080 3395 -2070
rect 3415 -2065 3425 -2060
rect 3740 -2060 3780 -2050
rect 3740 -2065 3750 -2060
rect 3415 -2080 3750 -2065
rect 3770 -2080 3780 -2060
rect -185 -2090 3780 -2080
rect -185 -2350 -165 -2090
rect -125 -2340 -60 -2330
rect -125 -2350 -115 -2340
rect -185 -2360 -115 -2350
rect -70 -2350 -60 -2340
rect 60 -2340 125 -2330
rect 60 -2350 70 -2340
rect -70 -2360 70 -2350
rect 115 -2350 125 -2340
rect 415 -2340 480 -2330
rect 415 -2350 425 -2340
rect 115 -2360 425 -2350
rect 470 -2350 480 -2340
rect 600 -2340 665 -2330
rect 600 -2350 610 -2340
rect 470 -2360 610 -2350
rect 655 -2350 665 -2340
rect 955 -2340 1020 -2330
rect 955 -2350 965 -2340
rect 655 -2360 965 -2350
rect 1010 -2350 1020 -2340
rect 1140 -2340 1205 -2330
rect 1140 -2350 1150 -2340
rect 1010 -2360 1150 -2350
rect 1195 -2350 1205 -2340
rect 1495 -2340 1560 -2330
rect 1495 -2350 1505 -2340
rect 1195 -2360 1505 -2350
rect 1550 -2350 1560 -2340
rect 1680 -2340 1745 -2330
rect 1680 -2350 1690 -2340
rect 1550 -2360 1690 -2350
rect 1735 -2350 1745 -2340
rect 2035 -2340 2100 -2330
rect 2035 -2350 2045 -2340
rect 1735 -2360 2045 -2350
rect 2090 -2350 2100 -2340
rect 2220 -2340 2285 -2330
rect 2220 -2350 2230 -2340
rect 2090 -2360 2230 -2350
rect 2275 -2350 2285 -2340
rect 2575 -2340 2640 -2330
rect 2575 -2350 2585 -2340
rect 2275 -2360 2585 -2350
rect 2630 -2350 2640 -2340
rect 2760 -2340 2825 -2330
rect 2760 -2350 2770 -2340
rect 2630 -2360 2770 -2350
rect 2815 -2350 2825 -2340
rect 3115 -2340 3180 -2330
rect 3115 -2350 3125 -2340
rect 2815 -2360 3125 -2350
rect 3170 -2350 3180 -2340
rect 3300 -2340 3365 -2330
rect 3300 -2350 3310 -2340
rect 3170 -2360 3310 -2350
rect 3355 -2350 3365 -2340
rect 3655 -2340 3720 -2330
rect 3655 -2350 3665 -2340
rect 3355 -2360 3665 -2350
rect 3710 -2360 3720 -2340
rect -185 -2370 3720 -2360
rect -185 -2425 3720 -2415
rect -185 -2435 -115 -2425
rect -185 -2665 -165 -2435
rect -125 -2445 -115 -2435
rect -70 -2435 70 -2425
rect -70 -2445 -60 -2435
rect -125 -2455 -60 -2445
rect 60 -2445 70 -2435
rect 115 -2435 425 -2425
rect 115 -2445 125 -2435
rect 60 -2455 125 -2445
rect 415 -2445 425 -2435
rect 470 -2435 610 -2425
rect 470 -2445 480 -2435
rect 415 -2455 480 -2445
rect 600 -2445 610 -2435
rect 655 -2435 965 -2425
rect 655 -2445 665 -2435
rect 600 -2455 665 -2445
rect 955 -2445 965 -2435
rect 1010 -2435 1150 -2425
rect 1010 -2445 1020 -2435
rect 955 -2455 1020 -2445
rect 1140 -2445 1150 -2435
rect 1195 -2435 1505 -2425
rect 1195 -2445 1205 -2435
rect 1140 -2455 1205 -2445
rect 1495 -2445 1505 -2435
rect 1550 -2435 1690 -2425
rect 1550 -2445 1560 -2435
rect 1495 -2455 1560 -2445
rect 1680 -2445 1690 -2435
rect 1735 -2435 2045 -2425
rect 1735 -2445 1745 -2435
rect 1680 -2455 1745 -2445
rect 2035 -2445 2045 -2435
rect 2090 -2435 2230 -2425
rect 2090 -2445 2100 -2435
rect 2035 -2455 2100 -2445
rect 2220 -2445 2230 -2435
rect 2275 -2435 2585 -2425
rect 2275 -2445 2285 -2435
rect 2220 -2455 2285 -2445
rect 2575 -2445 2585 -2435
rect 2630 -2435 2770 -2425
rect 2630 -2445 2640 -2435
rect 2575 -2455 2640 -2445
rect 2760 -2445 2770 -2435
rect 2815 -2435 3125 -2425
rect 2815 -2445 2825 -2435
rect 2760 -2455 2825 -2445
rect 3115 -2445 3125 -2435
rect 3170 -2435 3310 -2425
rect 3170 -2445 3180 -2435
rect 3115 -2455 3180 -2445
rect 3300 -2445 3310 -2435
rect 3355 -2435 3665 -2425
rect 3355 -2445 3365 -2435
rect 3300 -2455 3365 -2445
rect 3655 -2445 3665 -2435
rect 3710 -2445 3720 -2425
rect 3655 -2455 3720 -2445
rect 3760 -2665 3780 -2090
rect -185 -2675 3780 -2665
rect -185 -2695 -175 -2675
rect -155 -2685 155 -2675
rect -155 -2695 -145 -2685
rect -185 -2705 -145 -2695
rect 145 -2695 155 -2685
rect 175 -2685 365 -2675
rect 175 -2695 185 -2685
rect 145 -2705 185 -2695
rect 355 -2695 365 -2685
rect 385 -2685 695 -2675
rect 385 -2695 395 -2685
rect 355 -2705 395 -2695
rect 685 -2695 695 -2685
rect 715 -2685 905 -2675
rect 715 -2695 725 -2685
rect 685 -2705 725 -2695
rect 895 -2695 905 -2685
rect 925 -2685 1235 -2675
rect 925 -2695 935 -2685
rect 895 -2705 935 -2695
rect 1225 -2695 1235 -2685
rect 1255 -2685 1445 -2675
rect 1255 -2695 1265 -2685
rect 1225 -2705 1265 -2695
rect 1435 -2695 1445 -2685
rect 1465 -2685 1775 -2675
rect 1465 -2695 1475 -2685
rect 1435 -2705 1475 -2695
rect 1765 -2695 1775 -2685
rect 1795 -2685 1985 -2675
rect 1795 -2695 1805 -2685
rect 1765 -2705 1805 -2695
rect 1975 -2695 1985 -2685
rect 2005 -2685 2315 -2675
rect 2005 -2695 2015 -2685
rect 1975 -2705 2015 -2695
rect 2305 -2695 2315 -2685
rect 2335 -2685 2525 -2675
rect 2335 -2695 2345 -2685
rect 2305 -2705 2345 -2695
rect 2515 -2695 2525 -2685
rect 2545 -2685 2855 -2675
rect 2545 -2695 2555 -2685
rect 2515 -2705 2555 -2695
rect 2845 -2695 2855 -2685
rect 2875 -2685 3065 -2675
rect 2875 -2695 2885 -2685
rect 2845 -2705 2885 -2695
rect 3055 -2695 3065 -2685
rect 3085 -2685 3395 -2675
rect 3085 -2695 3095 -2685
rect 3055 -2705 3095 -2695
rect 3385 -2695 3395 -2685
rect 3415 -2685 3750 -2675
rect 3415 -2695 3425 -2685
rect 3385 -2705 3425 -2695
rect 3740 -2695 3750 -2685
rect 3770 -2695 3780 -2675
rect 3740 -2705 3780 -2695
rect -125 -2975 -60 -2965
rect -125 -2995 -115 -2975
rect -70 -2995 -60 -2975
rect -125 -3005 -60 -2995
rect 60 -2975 125 -2965
rect 60 -2995 70 -2975
rect 115 -2995 125 -2975
rect 415 -2975 480 -2965
rect 415 -2985 425 -2975
rect 60 -3005 125 -2995
rect 245 -2995 425 -2985
rect 470 -2995 480 -2975
rect 245 -3005 480 -2995
rect 600 -2975 665 -2965
rect 600 -2995 610 -2975
rect 655 -2995 665 -2975
rect 955 -2975 1020 -2965
rect 955 -2985 965 -2975
rect 600 -3005 665 -2995
rect 785 -2995 965 -2985
rect 1010 -2995 1020 -2975
rect 785 -3005 1020 -2995
rect 1140 -2975 1205 -2965
rect 1140 -2995 1150 -2975
rect 1195 -2995 1205 -2975
rect 1495 -2975 1560 -2965
rect 1495 -2985 1505 -2975
rect 1140 -3005 1205 -2995
rect 1325 -2995 1505 -2985
rect 1550 -2995 1560 -2975
rect 1325 -3005 1560 -2995
rect 1680 -2975 1745 -2965
rect 1680 -2995 1690 -2975
rect 1735 -2995 1745 -2975
rect 2035 -2975 2100 -2965
rect 2035 -2985 2045 -2975
rect 1680 -3005 1745 -2995
rect 1865 -2995 2045 -2985
rect 2090 -2995 2100 -2975
rect 1865 -3005 2100 -2995
rect 2220 -2975 2285 -2965
rect 2220 -2995 2230 -2975
rect 2275 -2995 2285 -2975
rect 2575 -2975 2640 -2965
rect 2575 -2985 2585 -2975
rect 2220 -3005 2285 -2995
rect 2405 -2995 2585 -2985
rect 2630 -2995 2640 -2975
rect 2405 -3005 2640 -2995
rect 2760 -2975 2825 -2965
rect 2760 -2995 2770 -2975
rect 2815 -2995 2825 -2975
rect 3115 -2975 3180 -2965
rect 3115 -2985 3125 -2975
rect 2760 -3005 2825 -2995
rect 2945 -2995 3125 -2985
rect 3170 -2995 3180 -2975
rect 2945 -3005 3180 -2995
rect 3300 -2975 3365 -2965
rect 3300 -2995 3310 -2975
rect 3355 -2995 3365 -2975
rect 3655 -2975 3720 -2965
rect 3655 -2985 3665 -2975
rect 3300 -3005 3365 -2995
rect 3470 -2995 3665 -2985
rect 3710 -2995 3720 -2975
rect 3470 -3005 3720 -2995
rect 145 -3260 185 -3250
rect -185 -3270 -145 -3260
rect -185 -3290 -175 -3270
rect -155 -3290 -145 -3270
rect 145 -3280 155 -3260
rect 175 -3280 185 -3260
rect 145 -3290 185 -3280
rect -185 -3300 -145 -3290
rect -185 -3810 -165 -3300
rect -125 -3525 -60 -3515
rect -125 -3545 -115 -3525
rect -70 -3545 -60 -3525
rect -125 -3555 -60 -3545
rect 60 -3525 125 -3515
rect 60 -3545 70 -3525
rect 115 -3545 125 -3525
rect 60 -3555 125 -3545
rect 165 -3800 185 -3290
rect 145 -3810 185 -3800
rect -185 -3820 -145 -3810
rect -185 -3840 -175 -3820
rect -155 -3840 -145 -3820
rect 145 -3830 155 -3810
rect 175 -3830 185 -3810
rect 145 -3840 185 -3830
rect -185 -3850 -145 -3840
rect -185 -4360 -165 -3850
rect -20 -3855 20 -3845
rect -20 -3925 -10 -3855
rect 10 -3925 20 -3855
rect -20 -3935 20 -3925
rect -125 -4075 -60 -4065
rect -125 -4095 -115 -4075
rect -70 -4095 -60 -4075
rect -125 -4105 -60 -4095
rect 60 -4075 125 -4065
rect 60 -4095 70 -4075
rect 115 -4095 125 -4075
rect 60 -4105 125 -4095
rect 165 -4350 185 -3840
rect 145 -4360 185 -4350
rect -185 -4370 -145 -4360
rect -185 -4390 -175 -4370
rect -155 -4390 -145 -4370
rect 145 -4380 155 -4360
rect 175 -4380 185 -4360
rect 145 -4390 185 -4380
rect -185 -4400 -145 -4390
rect -185 -4910 -165 -4400
rect -125 -4625 -60 -4615
rect -125 -4645 -115 -4625
rect -70 -4645 -60 -4625
rect -125 -4655 -60 -4645
rect 60 -4625 125 -4615
rect 60 -4645 70 -4625
rect 115 -4645 125 -4625
rect 60 -4655 125 -4645
rect 165 -4900 185 -4390
rect 145 -4910 185 -4900
rect -185 -4920 -145 -4910
rect -185 -4940 -175 -4920
rect -155 -4940 -145 -4920
rect 145 -4930 155 -4910
rect 175 -4930 185 -4910
rect 145 -4940 185 -4930
rect -185 -4950 -145 -4940
rect 245 -5165 265 -3005
rect 355 -3260 395 -3250
rect 355 -3280 365 -3260
rect 385 -3280 395 -3260
rect 355 -3290 395 -3280
rect 685 -3260 725 -3250
rect 685 -3280 695 -3260
rect 715 -3280 725 -3260
rect 685 -3290 725 -3280
rect 355 -3800 375 -3290
rect 415 -3525 480 -3515
rect 415 -3545 425 -3525
rect 470 -3545 480 -3525
rect 415 -3555 480 -3545
rect 600 -3525 665 -3515
rect 600 -3545 610 -3525
rect 655 -3545 665 -3525
rect 600 -3555 665 -3545
rect 705 -3800 725 -3290
rect 355 -3810 395 -3800
rect 355 -3830 365 -3810
rect 385 -3830 395 -3810
rect 355 -3840 395 -3830
rect 685 -3810 725 -3800
rect 685 -3830 695 -3810
rect 715 -3830 725 -3810
rect 685 -3840 725 -3830
rect 355 -4350 375 -3840
rect 520 -3855 560 -3845
rect 520 -3925 530 -3855
rect 550 -3925 560 -3855
rect 520 -3935 560 -3925
rect 415 -4075 480 -4065
rect 415 -4095 425 -4075
rect 470 -4095 480 -4075
rect 415 -4105 480 -4095
rect 600 -4075 665 -4065
rect 600 -4095 610 -4075
rect 655 -4095 665 -4075
rect 600 -4105 665 -4095
rect 705 -4350 725 -3840
rect 355 -4360 395 -4350
rect 355 -4380 365 -4360
rect 385 -4380 395 -4360
rect 355 -4390 395 -4380
rect 685 -4360 725 -4350
rect 685 -4380 695 -4360
rect 715 -4380 725 -4360
rect 685 -4390 725 -4380
rect 355 -4900 375 -4390
rect 415 -4625 480 -4615
rect 415 -4645 425 -4625
rect 470 -4645 480 -4625
rect 415 -4655 480 -4645
rect 600 -4625 665 -4615
rect 600 -4645 610 -4625
rect 655 -4645 665 -4625
rect 600 -4655 665 -4645
rect 705 -4900 725 -4390
rect 355 -4910 395 -4900
rect 355 -4930 365 -4910
rect 385 -4930 395 -4910
rect 355 -4940 395 -4930
rect 685 -4910 725 -4900
rect 685 -4930 695 -4910
rect 715 -4930 725 -4910
rect 685 -4940 725 -4930
rect 785 -5165 805 -3005
rect 895 -3260 935 -3250
rect 895 -3280 905 -3260
rect 925 -3280 935 -3260
rect 895 -3290 935 -3280
rect 1225 -3260 1265 -3250
rect 1225 -3280 1235 -3260
rect 1255 -3280 1265 -3260
rect 1225 -3290 1265 -3280
rect 895 -3800 915 -3290
rect 955 -3525 1020 -3515
rect 955 -3545 965 -3525
rect 1010 -3545 1020 -3525
rect 955 -3555 1020 -3545
rect 1140 -3525 1205 -3515
rect 1140 -3545 1150 -3525
rect 1195 -3545 1205 -3525
rect 1140 -3555 1205 -3545
rect 1245 -3800 1265 -3290
rect 895 -3810 935 -3800
rect 895 -3830 905 -3810
rect 925 -3830 935 -3810
rect 895 -3840 935 -3830
rect 1225 -3810 1265 -3800
rect 1225 -3830 1235 -3810
rect 1255 -3830 1265 -3810
rect 1225 -3840 1265 -3830
rect 895 -4350 915 -3840
rect 1060 -3855 1100 -3845
rect 1060 -3925 1070 -3855
rect 1090 -3925 1100 -3855
rect 1060 -3935 1100 -3925
rect 955 -4075 1020 -4065
rect 955 -4095 965 -4075
rect 1010 -4095 1020 -4075
rect 955 -4105 1020 -4095
rect 1140 -4075 1205 -4065
rect 1140 -4095 1150 -4075
rect 1195 -4095 1205 -4075
rect 1140 -4105 1205 -4095
rect 1245 -4350 1265 -3840
rect 895 -4360 935 -4350
rect 895 -4380 905 -4360
rect 925 -4380 935 -4360
rect 895 -4390 935 -4380
rect 1225 -4360 1265 -4350
rect 1225 -4380 1235 -4360
rect 1255 -4380 1265 -4360
rect 1225 -4390 1265 -4380
rect 895 -4900 915 -4390
rect 955 -4625 1020 -4615
rect 955 -4645 965 -4625
rect 1010 -4645 1020 -4625
rect 955 -4655 1020 -4645
rect 1140 -4625 1205 -4615
rect 1140 -4645 1150 -4625
rect 1195 -4645 1205 -4625
rect 1140 -4655 1205 -4645
rect 1245 -4900 1265 -4390
rect 895 -4910 935 -4900
rect 895 -4930 905 -4910
rect 925 -4930 935 -4910
rect 895 -4940 935 -4930
rect 1225 -4910 1265 -4900
rect 1225 -4930 1235 -4910
rect 1255 -4930 1265 -4910
rect 1225 -4940 1265 -4930
rect 1325 -5165 1345 -3005
rect 1435 -3260 1475 -3250
rect 1435 -3280 1445 -3260
rect 1465 -3280 1475 -3260
rect 1435 -3290 1475 -3280
rect 1765 -3260 1805 -3250
rect 1765 -3280 1775 -3260
rect 1795 -3280 1805 -3260
rect 1765 -3290 1805 -3280
rect 1435 -3800 1455 -3290
rect 1495 -3525 1560 -3515
rect 1495 -3545 1505 -3525
rect 1550 -3545 1560 -3525
rect 1495 -3555 1560 -3545
rect 1680 -3525 1745 -3515
rect 1680 -3545 1690 -3525
rect 1735 -3545 1745 -3525
rect 1680 -3555 1745 -3545
rect 1785 -3800 1805 -3290
rect 1435 -3810 1475 -3800
rect 1435 -3830 1445 -3810
rect 1465 -3830 1475 -3810
rect 1435 -3840 1475 -3830
rect 1765 -3810 1805 -3800
rect 1765 -3830 1775 -3810
rect 1795 -3830 1805 -3810
rect 1765 -3840 1805 -3830
rect 1435 -4350 1455 -3840
rect 1600 -3855 1640 -3845
rect 1600 -3925 1610 -3855
rect 1630 -3925 1640 -3855
rect 1600 -3935 1640 -3925
rect 1495 -4075 1560 -4065
rect 1495 -4095 1505 -4075
rect 1550 -4095 1560 -4075
rect 1495 -4105 1560 -4095
rect 1680 -4075 1745 -4065
rect 1680 -4095 1690 -4075
rect 1735 -4095 1745 -4075
rect 1680 -4105 1745 -4095
rect 1785 -4350 1805 -3840
rect 1435 -4360 1475 -4350
rect 1435 -4380 1445 -4360
rect 1465 -4380 1475 -4360
rect 1435 -4390 1475 -4380
rect 1765 -4360 1805 -4350
rect 1765 -4380 1775 -4360
rect 1795 -4380 1805 -4360
rect 1765 -4390 1805 -4380
rect 1435 -4900 1455 -4390
rect 1495 -4625 1560 -4615
rect 1495 -4645 1505 -4625
rect 1550 -4645 1560 -4625
rect 1495 -4655 1560 -4645
rect 1680 -4625 1745 -4615
rect 1680 -4645 1690 -4625
rect 1735 -4645 1745 -4625
rect 1680 -4655 1745 -4645
rect 1785 -4900 1805 -4390
rect 1435 -4910 1475 -4900
rect 1435 -4930 1445 -4910
rect 1465 -4930 1475 -4910
rect 1435 -4940 1475 -4930
rect 1765 -4910 1805 -4900
rect 1765 -4930 1775 -4910
rect 1795 -4930 1805 -4910
rect 1765 -4940 1805 -4930
rect 1865 -5165 1885 -3005
rect 1975 -3260 2015 -3250
rect 1975 -3280 1985 -3260
rect 2005 -3280 2015 -3260
rect 1975 -3290 2015 -3280
rect 2305 -3260 2345 -3250
rect 2305 -3280 2315 -3260
rect 2335 -3280 2345 -3260
rect 2305 -3290 2345 -3280
rect 1975 -3800 1995 -3290
rect 2035 -3525 2100 -3515
rect 2035 -3545 2045 -3525
rect 2090 -3545 2100 -3525
rect 2035 -3555 2100 -3545
rect 2220 -3525 2285 -3515
rect 2220 -3545 2230 -3525
rect 2275 -3545 2285 -3525
rect 2220 -3555 2285 -3545
rect 2325 -3800 2345 -3290
rect 1975 -3810 2015 -3800
rect 1975 -3830 1985 -3810
rect 2005 -3830 2015 -3810
rect 1975 -3840 2015 -3830
rect 2305 -3810 2345 -3800
rect 2305 -3830 2315 -3810
rect 2335 -3830 2345 -3810
rect 2305 -3840 2345 -3830
rect 1975 -4350 1995 -3840
rect 2140 -3855 2180 -3845
rect 2140 -3925 2150 -3855
rect 2170 -3925 2180 -3855
rect 2140 -3935 2180 -3925
rect 2035 -4075 2100 -4065
rect 2035 -4095 2045 -4075
rect 2090 -4095 2100 -4075
rect 2035 -4105 2100 -4095
rect 2220 -4075 2285 -4065
rect 2220 -4095 2230 -4075
rect 2275 -4095 2285 -4075
rect 2220 -4105 2285 -4095
rect 2325 -4350 2345 -3840
rect 1975 -4360 2015 -4350
rect 1975 -4380 1985 -4360
rect 2005 -4380 2015 -4360
rect 1975 -4390 2015 -4380
rect 2305 -4360 2345 -4350
rect 2305 -4380 2315 -4360
rect 2335 -4380 2345 -4360
rect 2305 -4390 2345 -4380
rect 1975 -4900 1995 -4390
rect 2035 -4625 2100 -4615
rect 2035 -4645 2045 -4625
rect 2090 -4645 2100 -4625
rect 2035 -4655 2100 -4645
rect 2220 -4625 2285 -4615
rect 2220 -4645 2230 -4625
rect 2275 -4645 2285 -4625
rect 2220 -4655 2285 -4645
rect 2325 -4900 2345 -4390
rect 1975 -4910 2015 -4900
rect 1975 -4930 1985 -4910
rect 2005 -4930 2015 -4910
rect 1975 -4940 2015 -4930
rect 2305 -4910 2345 -4900
rect 2305 -4930 2315 -4910
rect 2335 -4930 2345 -4910
rect 2305 -4940 2345 -4930
rect 2405 -5165 2425 -3005
rect 2515 -3260 2555 -3250
rect 2515 -3280 2525 -3260
rect 2545 -3280 2555 -3260
rect 2515 -3290 2555 -3280
rect 2845 -3260 2885 -3250
rect 2845 -3280 2855 -3260
rect 2875 -3280 2885 -3260
rect 2845 -3290 2885 -3280
rect 2515 -3800 2535 -3290
rect 2575 -3525 2640 -3515
rect 2575 -3545 2585 -3525
rect 2630 -3545 2640 -3525
rect 2575 -3555 2640 -3545
rect 2760 -3525 2825 -3515
rect 2760 -3545 2770 -3525
rect 2815 -3545 2825 -3525
rect 2760 -3555 2825 -3545
rect 2865 -3800 2885 -3290
rect 2515 -3810 2555 -3800
rect 2515 -3830 2525 -3810
rect 2545 -3830 2555 -3810
rect 2515 -3840 2555 -3830
rect 2845 -3810 2885 -3800
rect 2845 -3830 2855 -3810
rect 2875 -3830 2885 -3810
rect 2845 -3840 2885 -3830
rect 2515 -4350 2535 -3840
rect 2680 -3855 2720 -3845
rect 2680 -3925 2690 -3855
rect 2710 -3925 2720 -3855
rect 2680 -3935 2720 -3925
rect 2575 -4075 2640 -4065
rect 2575 -4095 2585 -4075
rect 2630 -4095 2640 -4075
rect 2575 -4105 2640 -4095
rect 2760 -4075 2825 -4065
rect 2760 -4095 2770 -4075
rect 2815 -4095 2825 -4075
rect 2760 -4105 2825 -4095
rect 2865 -4350 2885 -3840
rect 2515 -4360 2555 -4350
rect 2515 -4380 2525 -4360
rect 2545 -4380 2555 -4360
rect 2515 -4390 2555 -4380
rect 2845 -4360 2885 -4350
rect 2845 -4380 2855 -4360
rect 2875 -4380 2885 -4360
rect 2845 -4390 2885 -4380
rect 2515 -4900 2535 -4390
rect 2575 -4625 2640 -4615
rect 2575 -4645 2585 -4625
rect 2630 -4645 2640 -4625
rect 2575 -4655 2640 -4645
rect 2760 -4625 2825 -4615
rect 2760 -4645 2770 -4625
rect 2815 -4645 2825 -4625
rect 2760 -4655 2825 -4645
rect 2865 -4900 2885 -4390
rect 2515 -4910 2555 -4900
rect 2515 -4930 2525 -4910
rect 2545 -4930 2555 -4910
rect 2515 -4940 2555 -4930
rect 2845 -4910 2885 -4900
rect 2845 -4930 2855 -4910
rect 2875 -4930 2885 -4910
rect 2845 -4940 2885 -4930
rect 2945 -5165 2965 -3005
rect 3055 -3260 3095 -3250
rect 3055 -3280 3065 -3260
rect 3085 -3280 3095 -3260
rect 3055 -3290 3095 -3280
rect 3385 -3260 3425 -3250
rect 3385 -3280 3395 -3260
rect 3415 -3280 3425 -3260
rect 3385 -3290 3425 -3280
rect 3055 -3800 3075 -3290
rect 3115 -3525 3180 -3515
rect 3115 -3545 3125 -3525
rect 3170 -3545 3180 -3525
rect 3115 -3555 3180 -3545
rect 3300 -3525 3365 -3515
rect 3300 -3545 3310 -3525
rect 3355 -3545 3365 -3525
rect 3300 -3555 3365 -3545
rect 3405 -3800 3425 -3290
rect 3055 -3810 3095 -3800
rect 3055 -3830 3065 -3810
rect 3085 -3830 3095 -3810
rect 3055 -3840 3095 -3830
rect 3385 -3810 3425 -3800
rect 3385 -3830 3395 -3810
rect 3415 -3830 3425 -3810
rect 3385 -3840 3425 -3830
rect 3055 -4350 3075 -3840
rect 3220 -3855 3260 -3845
rect 3220 -3925 3230 -3855
rect 3250 -3925 3260 -3855
rect 3220 -3935 3260 -3925
rect 3115 -4075 3180 -4065
rect 3115 -4095 3125 -4075
rect 3170 -4095 3180 -4075
rect 3115 -4105 3180 -4095
rect 3300 -4075 3365 -4065
rect 3300 -4095 3310 -4075
rect 3355 -4095 3365 -4075
rect 3300 -4105 3365 -4095
rect 3405 -4350 3425 -3840
rect 3055 -4360 3095 -4350
rect 3055 -4380 3065 -4360
rect 3085 -4380 3095 -4360
rect 3055 -4390 3095 -4380
rect 3385 -4360 3425 -4350
rect 3385 -4380 3395 -4360
rect 3415 -4380 3425 -4360
rect 3385 -4390 3425 -4380
rect 3055 -4900 3075 -4390
rect 3115 -4625 3180 -4615
rect 3115 -4645 3125 -4625
rect 3170 -4645 3180 -4625
rect 3115 -4655 3180 -4645
rect 3300 -4625 3365 -4615
rect 3300 -4645 3310 -4625
rect 3355 -4645 3365 -4625
rect 3300 -4655 3365 -4645
rect 3405 -4900 3425 -4390
rect 3055 -4910 3095 -4900
rect 3055 -4930 3065 -4910
rect 3085 -4930 3095 -4910
rect 3055 -4940 3095 -4930
rect 3385 -4910 3425 -4900
rect 3385 -4930 3395 -4910
rect 3415 -4930 3425 -4910
rect 3385 -4940 3425 -4930
rect -125 -5175 -60 -5165
rect -125 -5195 -115 -5175
rect -70 -5195 -60 -5175
rect -125 -5205 -60 -5195
rect 60 -5175 265 -5165
rect 60 -5195 70 -5175
rect 115 -5185 265 -5175
rect 415 -5175 480 -5165
rect 115 -5195 125 -5185
rect 60 -5205 125 -5195
rect 415 -5195 425 -5175
rect 470 -5195 480 -5175
rect 415 -5205 480 -5195
rect 600 -5175 805 -5165
rect 600 -5195 610 -5175
rect 655 -5185 805 -5175
rect 955 -5175 1020 -5165
rect 655 -5195 665 -5185
rect 600 -5205 665 -5195
rect 955 -5195 965 -5175
rect 1010 -5195 1020 -5175
rect 955 -5205 1020 -5195
rect 1140 -5175 1345 -5165
rect 1140 -5195 1150 -5175
rect 1195 -5185 1345 -5175
rect 1495 -5175 1560 -5165
rect 1195 -5195 1205 -5185
rect 1140 -5205 1205 -5195
rect 1495 -5195 1505 -5175
rect 1550 -5195 1560 -5175
rect 1495 -5205 1560 -5195
rect 1680 -5175 1885 -5165
rect 1680 -5195 1690 -5175
rect 1735 -5185 1885 -5175
rect 2035 -5175 2100 -5165
rect 1735 -5195 1745 -5185
rect 1680 -5205 1745 -5195
rect 2035 -5195 2045 -5175
rect 2090 -5195 2100 -5175
rect 2035 -5205 2100 -5195
rect 2220 -5175 2425 -5165
rect 2220 -5195 2230 -5175
rect 2275 -5185 2425 -5175
rect 2575 -5175 2640 -5165
rect 2275 -5195 2285 -5185
rect 2220 -5205 2285 -5195
rect 2575 -5195 2585 -5175
rect 2630 -5195 2640 -5175
rect 2575 -5205 2640 -5195
rect 2760 -5175 2965 -5165
rect 2760 -5195 2770 -5175
rect 2815 -5185 2965 -5175
rect 3115 -5175 3180 -5165
rect 2815 -5195 2825 -5185
rect 2760 -5205 2825 -5195
rect 3115 -5195 3125 -5175
rect 3170 -5195 3180 -5175
rect 3115 -5205 3180 -5195
rect 3300 -5175 3365 -5165
rect 3300 -5195 3310 -5175
rect 3355 -5185 3365 -5175
rect 3470 -5185 3490 -3005
rect 3740 -3260 3780 -3250
rect 3740 -3280 3750 -3260
rect 3770 -3280 3780 -3260
rect 3740 -3290 3780 -3280
rect 3655 -3525 3720 -3515
rect 3655 -3545 3665 -3525
rect 3710 -3545 3720 -3525
rect 3655 -3555 3720 -3545
rect 3760 -3800 3780 -3290
rect 3740 -3810 3780 -3800
rect 3740 -3830 3750 -3810
rect 3770 -3830 3780 -3810
rect 3740 -3840 3780 -3830
rect 3655 -4075 3720 -4065
rect 3655 -4095 3665 -4075
rect 3710 -4095 3720 -4075
rect 3655 -4105 3720 -4095
rect 3760 -4350 3780 -3840
rect 3740 -4360 3780 -4350
rect 3740 -4380 3750 -4360
rect 3770 -4380 3780 -4360
rect 3740 -4390 3780 -4380
rect 3655 -4625 3720 -4615
rect 3655 -4645 3665 -4625
rect 3710 -4645 3720 -4625
rect 3655 -4655 3720 -4645
rect 3760 -4900 3780 -4390
rect 3740 -4910 3780 -4900
rect 3740 -4930 3750 -4910
rect 3770 -4930 3780 -4910
rect 3740 -4940 3780 -4930
rect 3355 -5195 3490 -5185
rect 3300 -5205 3490 -5195
rect 3655 -5175 3720 -5165
rect 3655 -5195 3665 -5175
rect 3710 -5195 3720 -5175
rect 3655 -5205 3720 -5195
rect -125 -5275 -105 -5205
rect 415 -5275 435 -5205
rect 955 -5275 975 -5205
rect 1495 -5275 1515 -5205
rect 2035 -5275 2055 -5205
rect 2575 -5275 2595 -5205
rect 3115 -5275 3135 -5205
rect -125 -5295 80 -5275
rect -125 -5320 -105 -5295
rect 60 -5320 80 -5295
rect 415 -5295 620 -5275
rect 415 -5320 435 -5295
rect 600 -5320 620 -5295
rect 955 -5295 1160 -5275
rect 955 -5320 975 -5295
rect 1140 -5320 1160 -5295
rect 1495 -5295 1700 -5275
rect 1495 -5320 1515 -5295
rect 1680 -5320 1700 -5295
rect 2035 -5295 2240 -5275
rect 2035 -5320 2055 -5295
rect 2220 -5320 2240 -5295
rect 2575 -5295 2780 -5275
rect 2575 -5320 2595 -5295
rect 2760 -5320 2780 -5295
rect 3115 -5295 3320 -5275
rect 3115 -5320 3135 -5295
rect 3300 -5320 3320 -5295
rect -125 -5330 -60 -5320
rect -125 -5350 -115 -5330
rect -70 -5350 -60 -5330
rect -125 -5360 -60 -5350
rect 60 -5330 125 -5320
rect 60 -5350 70 -5330
rect 115 -5350 125 -5330
rect 60 -5360 125 -5350
rect 415 -5330 480 -5320
rect 415 -5350 425 -5330
rect 470 -5350 480 -5330
rect 415 -5360 480 -5350
rect 600 -5330 665 -5320
rect 600 -5350 610 -5330
rect 655 -5350 665 -5330
rect 600 -5360 665 -5350
rect 955 -5330 1020 -5320
rect 955 -5350 965 -5330
rect 1010 -5350 1020 -5330
rect 955 -5360 1020 -5350
rect 1140 -5330 1205 -5320
rect 1140 -5350 1150 -5330
rect 1195 -5350 1205 -5330
rect 1140 -5360 1205 -5350
rect 1495 -5330 1560 -5320
rect 1495 -5350 1505 -5330
rect 1550 -5350 1560 -5330
rect 1495 -5360 1560 -5350
rect 1680 -5330 1745 -5320
rect 1680 -5350 1690 -5330
rect 1735 -5350 1745 -5330
rect 1680 -5360 1745 -5350
rect 2035 -5330 2100 -5320
rect 2035 -5350 2045 -5330
rect 2090 -5350 2100 -5330
rect 2035 -5360 2100 -5350
rect 2220 -5330 2285 -5320
rect 2220 -5350 2230 -5330
rect 2275 -5350 2285 -5330
rect 2220 -5360 2285 -5350
rect 2575 -5330 2640 -5320
rect 2575 -5350 2585 -5330
rect 2630 -5350 2640 -5330
rect 2575 -5360 2640 -5350
rect 2760 -5330 2825 -5320
rect 2760 -5350 2770 -5330
rect 2815 -5350 2825 -5330
rect 2760 -5360 2825 -5350
rect 3115 -5330 3180 -5320
rect 3115 -5350 3125 -5330
rect 3170 -5350 3180 -5330
rect 3115 -5360 3180 -5350
rect 3300 -5330 3365 -5320
rect 3300 -5350 3310 -5330
rect 3355 -5350 3365 -5330
rect 3300 -5360 3365 -5350
rect -185 -5620 -145 -5610
rect -185 -5640 -175 -5620
rect -155 -5640 -145 -5620
rect -185 -5650 -145 -5640
rect 145 -5620 185 -5610
rect 145 -5640 155 -5620
rect 175 -5640 185 -5620
rect 145 -5650 185 -5640
rect -185 -6160 -165 -5650
rect -125 -5880 -60 -5870
rect -125 -5900 -115 -5880
rect -70 -5900 -60 -5880
rect -125 -5910 -60 -5900
rect 60 -5880 125 -5870
rect 60 -5900 70 -5880
rect 115 -5900 125 -5880
rect 60 -5910 125 -5900
rect 165 -6160 185 -5650
rect -185 -6170 -145 -6160
rect -185 -6190 -175 -6170
rect -155 -6190 -145 -6170
rect -185 -6200 -145 -6190
rect 145 -6170 185 -6160
rect 145 -6190 155 -6170
rect 175 -6190 185 -6170
rect 145 -6200 185 -6190
rect -185 -6710 -165 -6200
rect -125 -6430 -60 -6420
rect -125 -6450 -115 -6430
rect -70 -6450 -60 -6430
rect -125 -6460 -60 -6450
rect 60 -6430 125 -6420
rect 60 -6450 70 -6430
rect 115 -6450 125 -6430
rect 60 -6460 125 -6450
rect 165 -6710 185 -6200
rect -185 -6720 -145 -6710
rect -185 -6740 -175 -6720
rect -155 -6740 -145 -6720
rect -185 -6750 -145 -6740
rect 145 -6720 185 -6710
rect 145 -6740 155 -6720
rect 175 -6740 185 -6720
rect 145 -6750 185 -6740
rect -185 -7260 -165 -6750
rect -20 -6760 20 -6750
rect -20 -6830 -10 -6760
rect 10 -6830 20 -6760
rect -20 -6840 20 -6830
rect -125 -6980 -60 -6970
rect -125 -7000 -115 -6980
rect -70 -7000 -60 -6980
rect -125 -7010 -60 -7000
rect 60 -6980 125 -6970
rect 60 -7000 70 -6980
rect 115 -7000 125 -6980
rect 60 -7010 125 -7000
rect 165 -7135 185 -6750
rect 355 -5620 395 -5610
rect 355 -5640 365 -5620
rect 385 -5640 395 -5620
rect 355 -5650 395 -5640
rect 685 -5620 725 -5610
rect 685 -5640 695 -5620
rect 715 -5640 725 -5620
rect 685 -5650 725 -5640
rect 355 -6160 375 -5650
rect 415 -5880 480 -5870
rect 415 -5900 425 -5880
rect 470 -5900 480 -5880
rect 415 -5910 480 -5900
rect 600 -5880 665 -5870
rect 600 -5900 610 -5880
rect 655 -5900 665 -5880
rect 600 -5910 665 -5900
rect 705 -6160 725 -5650
rect 355 -6170 395 -6160
rect 355 -6190 365 -6170
rect 385 -6190 395 -6170
rect 355 -6200 395 -6190
rect 685 -6170 725 -6160
rect 685 -6190 695 -6170
rect 715 -6190 725 -6170
rect 685 -6200 725 -6190
rect 355 -6710 375 -6200
rect 415 -6430 480 -6420
rect 415 -6450 425 -6430
rect 470 -6450 480 -6430
rect 415 -6460 480 -6450
rect 600 -6430 665 -6420
rect 600 -6450 610 -6430
rect 655 -6450 665 -6430
rect 600 -6460 665 -6450
rect 705 -6710 725 -6200
rect 355 -6720 395 -6710
rect 355 -6740 365 -6720
rect 385 -6740 395 -6720
rect 355 -6750 395 -6740
rect 685 -6720 725 -6710
rect 685 -6740 695 -6720
rect 715 -6740 725 -6720
rect 685 -6750 725 -6740
rect 355 -7060 375 -6750
rect 520 -6760 560 -6750
rect 520 -6830 530 -6760
rect 550 -6830 560 -6760
rect 520 -6840 560 -6830
rect 415 -6980 480 -6970
rect 415 -7000 425 -6980
rect 470 -7000 480 -6980
rect 415 -7010 480 -7000
rect 600 -6980 665 -6970
rect 600 -7000 610 -6980
rect 655 -7000 665 -6980
rect 600 -7010 665 -7000
rect 280 -7070 375 -7060
rect 280 -7100 290 -7070
rect 345 -7100 375 -7070
rect 280 -7110 375 -7100
rect 165 -7145 260 -7135
rect 165 -7175 195 -7145
rect 250 -7175 260 -7145
rect 165 -7185 260 -7175
rect 165 -7260 185 -7185
rect -185 -7270 -145 -7260
rect -185 -7290 -175 -7270
rect -155 -7290 -145 -7270
rect -185 -7300 -145 -7290
rect 145 -7270 185 -7260
rect 145 -7290 155 -7270
rect 175 -7290 185 -7270
rect 145 -7300 185 -7290
rect 355 -7260 375 -7110
rect 705 -7135 725 -6750
rect 895 -5620 935 -5610
rect 895 -5640 905 -5620
rect 925 -5640 935 -5620
rect 895 -5650 935 -5640
rect 1225 -5620 1265 -5610
rect 1225 -5640 1235 -5620
rect 1255 -5640 1265 -5620
rect 1225 -5650 1265 -5640
rect 895 -6160 915 -5650
rect 955 -5880 1020 -5870
rect 955 -5900 965 -5880
rect 1010 -5900 1020 -5880
rect 955 -5910 1020 -5900
rect 1140 -5880 1205 -5870
rect 1140 -5900 1150 -5880
rect 1195 -5900 1205 -5880
rect 1140 -5910 1205 -5900
rect 1245 -6160 1265 -5650
rect 895 -6170 935 -6160
rect 895 -6190 905 -6170
rect 925 -6190 935 -6170
rect 895 -6200 935 -6190
rect 1225 -6170 1265 -6160
rect 1225 -6190 1235 -6170
rect 1255 -6190 1265 -6170
rect 1225 -6200 1265 -6190
rect 895 -6710 915 -6200
rect 955 -6430 1020 -6420
rect 955 -6450 965 -6430
rect 1010 -6450 1020 -6430
rect 955 -6460 1020 -6450
rect 1140 -6430 1205 -6420
rect 1140 -6450 1150 -6430
rect 1195 -6450 1205 -6430
rect 1140 -6460 1205 -6450
rect 1245 -6710 1265 -6200
rect 895 -6720 935 -6710
rect 895 -6740 905 -6720
rect 925 -6740 935 -6720
rect 895 -6750 935 -6740
rect 1225 -6720 1265 -6710
rect 1225 -6740 1235 -6720
rect 1255 -6740 1265 -6720
rect 1225 -6750 1265 -6740
rect 895 -7060 915 -6750
rect 1060 -6760 1100 -6750
rect 1060 -6830 1070 -6760
rect 1090 -6830 1100 -6760
rect 1060 -6840 1100 -6830
rect 955 -6980 1020 -6970
rect 955 -7000 965 -6980
rect 1010 -7000 1020 -6980
rect 955 -7010 1020 -7000
rect 1140 -6980 1205 -6970
rect 1140 -7000 1150 -6980
rect 1195 -7000 1205 -6980
rect 1140 -7010 1205 -7000
rect 820 -7070 915 -7060
rect 820 -7100 830 -7070
rect 885 -7100 915 -7070
rect 820 -7110 915 -7100
rect 705 -7145 800 -7135
rect 705 -7175 735 -7145
rect 790 -7175 800 -7145
rect 705 -7185 800 -7175
rect 705 -7260 725 -7185
rect 355 -7270 395 -7260
rect 355 -7290 365 -7270
rect 385 -7290 395 -7270
rect 355 -7300 395 -7290
rect 685 -7270 725 -7260
rect 685 -7290 695 -7270
rect 715 -7290 725 -7270
rect 685 -7300 725 -7290
rect 895 -7260 915 -7110
rect 1245 -7135 1265 -6750
rect 1435 -5620 1475 -5610
rect 1435 -5640 1445 -5620
rect 1465 -5640 1475 -5620
rect 1435 -5650 1475 -5640
rect 1765 -5620 1805 -5610
rect 1765 -5640 1775 -5620
rect 1795 -5640 1805 -5620
rect 1765 -5650 1805 -5640
rect 1435 -6160 1455 -5650
rect 1495 -5880 1560 -5870
rect 1495 -5900 1505 -5880
rect 1550 -5900 1560 -5880
rect 1495 -5910 1560 -5900
rect 1680 -5880 1745 -5870
rect 1680 -5900 1690 -5880
rect 1735 -5900 1745 -5880
rect 1680 -5910 1745 -5900
rect 1785 -6160 1805 -5650
rect 1435 -6170 1475 -6160
rect 1435 -6190 1445 -6170
rect 1465 -6190 1475 -6170
rect 1435 -6200 1475 -6190
rect 1765 -6170 1805 -6160
rect 1765 -6190 1775 -6170
rect 1795 -6190 1805 -6170
rect 1765 -6200 1805 -6190
rect 1435 -6710 1455 -6200
rect 1495 -6430 1560 -6420
rect 1495 -6450 1505 -6430
rect 1550 -6450 1560 -6430
rect 1495 -6460 1560 -6450
rect 1680 -6430 1745 -6420
rect 1680 -6450 1690 -6430
rect 1735 -6450 1745 -6430
rect 1680 -6460 1745 -6450
rect 1785 -6710 1805 -6200
rect 1435 -6720 1475 -6710
rect 1435 -6740 1445 -6720
rect 1465 -6740 1475 -6720
rect 1435 -6750 1475 -6740
rect 1765 -6720 1805 -6710
rect 1765 -6740 1775 -6720
rect 1795 -6740 1805 -6720
rect 1765 -6750 1805 -6740
rect 1435 -7060 1455 -6750
rect 1600 -6760 1640 -6750
rect 1600 -6830 1610 -6760
rect 1630 -6830 1640 -6760
rect 1600 -6840 1640 -6830
rect 1495 -6980 1560 -6970
rect 1495 -7000 1505 -6980
rect 1550 -7000 1560 -6980
rect 1495 -7010 1560 -7000
rect 1680 -6980 1745 -6970
rect 1680 -7000 1690 -6980
rect 1735 -7000 1745 -6980
rect 1680 -7010 1745 -7000
rect 1360 -7070 1455 -7060
rect 1360 -7100 1370 -7070
rect 1425 -7100 1455 -7070
rect 1360 -7110 1455 -7100
rect 1245 -7145 1340 -7135
rect 1245 -7175 1275 -7145
rect 1330 -7175 1340 -7145
rect 1245 -7185 1340 -7175
rect 1245 -7260 1265 -7185
rect 895 -7270 935 -7260
rect 895 -7290 905 -7270
rect 925 -7290 935 -7270
rect 895 -7300 935 -7290
rect 1225 -7270 1265 -7260
rect 1225 -7290 1235 -7270
rect 1255 -7290 1265 -7270
rect 1225 -7300 1265 -7290
rect 1435 -7260 1455 -7110
rect 1785 -7135 1805 -6750
rect 1975 -5620 2015 -5610
rect 1975 -5640 1985 -5620
rect 2005 -5640 2015 -5620
rect 1975 -5650 2015 -5640
rect 2305 -5620 2345 -5610
rect 2305 -5640 2315 -5620
rect 2335 -5640 2345 -5620
rect 2305 -5650 2345 -5640
rect 1975 -6160 1995 -5650
rect 2035 -5880 2100 -5870
rect 2035 -5900 2045 -5880
rect 2090 -5900 2100 -5880
rect 2035 -5910 2100 -5900
rect 2220 -5880 2285 -5870
rect 2220 -5900 2230 -5880
rect 2275 -5900 2285 -5880
rect 2220 -5910 2285 -5900
rect 2325 -6160 2345 -5650
rect 1975 -6170 2015 -6160
rect 1975 -6190 1985 -6170
rect 2005 -6190 2015 -6170
rect 1975 -6200 2015 -6190
rect 2305 -6170 2345 -6160
rect 2305 -6190 2315 -6170
rect 2335 -6190 2345 -6170
rect 2305 -6200 2345 -6190
rect 1975 -6710 1995 -6200
rect 2035 -6430 2100 -6420
rect 2035 -6450 2045 -6430
rect 2090 -6450 2100 -6430
rect 2035 -6460 2100 -6450
rect 2220 -6430 2285 -6420
rect 2220 -6450 2230 -6430
rect 2275 -6450 2285 -6430
rect 2220 -6460 2285 -6450
rect 2325 -6710 2345 -6200
rect 1975 -6720 2015 -6710
rect 1975 -6740 1985 -6720
rect 2005 -6740 2015 -6720
rect 1975 -6750 2015 -6740
rect 2305 -6720 2345 -6710
rect 2305 -6740 2315 -6720
rect 2335 -6740 2345 -6720
rect 2305 -6750 2345 -6740
rect 1975 -7060 1995 -6750
rect 2140 -6760 2180 -6750
rect 2140 -6830 2150 -6760
rect 2170 -6830 2180 -6760
rect 2140 -6840 2180 -6830
rect 2035 -6980 2100 -6970
rect 2035 -7000 2045 -6980
rect 2090 -7000 2100 -6980
rect 2035 -7010 2100 -7000
rect 2220 -6980 2285 -6970
rect 2220 -7000 2230 -6980
rect 2275 -7000 2285 -6980
rect 2220 -7010 2285 -7000
rect 1900 -7070 1995 -7060
rect 1900 -7100 1910 -7070
rect 1965 -7100 1995 -7070
rect 1900 -7110 1995 -7100
rect 1785 -7145 1880 -7135
rect 1785 -7175 1815 -7145
rect 1870 -7175 1880 -7145
rect 1785 -7185 1880 -7175
rect 1785 -7260 1805 -7185
rect 1435 -7270 1475 -7260
rect 1435 -7290 1445 -7270
rect 1465 -7290 1475 -7270
rect 1435 -7300 1475 -7290
rect 1765 -7270 1805 -7260
rect 1765 -7290 1775 -7270
rect 1795 -7290 1805 -7270
rect 1765 -7300 1805 -7290
rect 1975 -7260 1995 -7110
rect 2325 -7135 2345 -6750
rect 2515 -5620 2555 -5610
rect 2515 -5640 2525 -5620
rect 2545 -5640 2555 -5620
rect 2515 -5650 2555 -5640
rect 2845 -5620 2885 -5610
rect 2845 -5640 2855 -5620
rect 2875 -5640 2885 -5620
rect 2845 -5650 2885 -5640
rect 2515 -6160 2535 -5650
rect 2575 -5880 2640 -5870
rect 2575 -5900 2585 -5880
rect 2630 -5900 2640 -5880
rect 2575 -5910 2640 -5900
rect 2760 -5880 2825 -5870
rect 2760 -5900 2770 -5880
rect 2815 -5900 2825 -5880
rect 2760 -5910 2825 -5900
rect 2865 -6160 2885 -5650
rect 2515 -6170 2555 -6160
rect 2515 -6190 2525 -6170
rect 2545 -6190 2555 -6170
rect 2515 -6200 2555 -6190
rect 2845 -6170 2885 -6160
rect 2845 -6190 2855 -6170
rect 2875 -6190 2885 -6170
rect 2845 -6200 2885 -6190
rect 2515 -6710 2535 -6200
rect 2575 -6430 2640 -6420
rect 2575 -6450 2585 -6430
rect 2630 -6450 2640 -6430
rect 2575 -6460 2640 -6450
rect 2760 -6430 2825 -6420
rect 2760 -6450 2770 -6430
rect 2815 -6450 2825 -6430
rect 2760 -6460 2825 -6450
rect 2865 -6710 2885 -6200
rect 2515 -6720 2555 -6710
rect 2515 -6740 2525 -6720
rect 2545 -6740 2555 -6720
rect 2515 -6750 2555 -6740
rect 2845 -6720 2885 -6710
rect 2845 -6740 2855 -6720
rect 2875 -6740 2885 -6720
rect 2845 -6750 2885 -6740
rect 2515 -7060 2535 -6750
rect 2680 -6760 2720 -6750
rect 2680 -6830 2690 -6760
rect 2710 -6830 2720 -6760
rect 2680 -6840 2720 -6830
rect 2575 -6980 2640 -6970
rect 2575 -7000 2585 -6980
rect 2630 -7000 2640 -6980
rect 2575 -7010 2640 -7000
rect 2760 -6980 2825 -6970
rect 2760 -7000 2770 -6980
rect 2815 -7000 2825 -6980
rect 2760 -7010 2825 -7000
rect 2440 -7070 2535 -7060
rect 2440 -7100 2450 -7070
rect 2505 -7100 2535 -7070
rect 2440 -7110 2535 -7100
rect 2325 -7145 2420 -7135
rect 2325 -7175 2355 -7145
rect 2410 -7175 2420 -7145
rect 2325 -7185 2420 -7175
rect 2325 -7260 2345 -7185
rect 1975 -7270 2015 -7260
rect 1975 -7290 1985 -7270
rect 2005 -7290 2015 -7270
rect 1975 -7300 2015 -7290
rect 2305 -7270 2345 -7260
rect 2305 -7290 2315 -7270
rect 2335 -7290 2345 -7270
rect 2305 -7300 2345 -7290
rect 2515 -7260 2535 -7110
rect 2865 -7135 2885 -6750
rect 3055 -5620 3095 -5610
rect 3055 -5640 3065 -5620
rect 3085 -5640 3095 -5620
rect 3055 -5650 3095 -5640
rect 3385 -5620 3425 -5610
rect 3385 -5640 3395 -5620
rect 3415 -5640 3425 -5620
rect 3385 -5650 3425 -5640
rect 3055 -6160 3075 -5650
rect 3115 -5880 3180 -5870
rect 3115 -5900 3125 -5880
rect 3170 -5900 3180 -5880
rect 3115 -5910 3180 -5900
rect 3300 -5880 3365 -5870
rect 3300 -5900 3310 -5880
rect 3355 -5900 3365 -5880
rect 3300 -5910 3365 -5900
rect 3405 -6160 3425 -5650
rect 3055 -6170 3095 -6160
rect 3055 -6190 3065 -6170
rect 3085 -6190 3095 -6170
rect 3055 -6200 3095 -6190
rect 3385 -6170 3425 -6160
rect 3385 -6190 3395 -6170
rect 3415 -6190 3425 -6170
rect 3385 -6200 3425 -6190
rect 3055 -6710 3075 -6200
rect 3115 -6430 3180 -6420
rect 3115 -6450 3125 -6430
rect 3170 -6450 3180 -6430
rect 3115 -6460 3180 -6450
rect 3300 -6430 3365 -6420
rect 3300 -6450 3310 -6430
rect 3355 -6450 3365 -6430
rect 3300 -6460 3365 -6450
rect 3405 -6710 3425 -6200
rect 3055 -6720 3095 -6710
rect 3055 -6740 3065 -6720
rect 3085 -6740 3095 -6720
rect 3055 -6750 3095 -6740
rect 3385 -6720 3425 -6710
rect 3385 -6740 3395 -6720
rect 3415 -6740 3425 -6720
rect 3385 -6750 3425 -6740
rect 3055 -7060 3075 -6750
rect 3220 -6760 3260 -6750
rect 3220 -6830 3230 -6760
rect 3250 -6830 3260 -6760
rect 3220 -6840 3260 -6830
rect 3115 -6980 3180 -6970
rect 3115 -7000 3125 -6980
rect 3170 -7000 3180 -6980
rect 3115 -7010 3180 -7000
rect 3300 -6980 3365 -6970
rect 3300 -7000 3310 -6980
rect 3355 -7000 3365 -6980
rect 3300 -7010 3365 -7000
rect 2980 -7070 3075 -7060
rect 2980 -7100 2990 -7070
rect 3045 -7100 3075 -7070
rect 2980 -7110 3075 -7100
rect 2865 -7145 2960 -7135
rect 2865 -7175 2895 -7145
rect 2950 -7175 2960 -7145
rect 2865 -7185 2960 -7175
rect 2865 -7260 2885 -7185
rect 2515 -7270 2555 -7260
rect 2515 -7290 2525 -7270
rect 2545 -7290 2555 -7270
rect 2515 -7300 2555 -7290
rect 2845 -7270 2885 -7260
rect 2845 -7290 2855 -7270
rect 2875 -7290 2885 -7270
rect 2845 -7300 2885 -7290
rect 3055 -7260 3075 -7110
rect 3405 -7060 3425 -6750
rect 3405 -7070 3500 -7060
rect 3405 -7100 3435 -7070
rect 3490 -7100 3500 -7070
rect 3405 -7110 3500 -7100
rect 3405 -7260 3425 -7110
rect 3055 -7270 3095 -7260
rect 3055 -7290 3065 -7270
rect 3085 -7290 3095 -7270
rect 3055 -7300 3095 -7290
rect 3385 -7270 3425 -7260
rect 3385 -7290 3395 -7270
rect 3415 -7290 3425 -7270
rect 3385 -7300 3425 -7290
rect -125 -7530 -60 -7520
rect -125 -7550 -115 -7530
rect -70 -7550 -60 -7530
rect -125 -7560 -60 -7550
rect 60 -7530 125 -7520
rect 60 -7550 70 -7530
rect 115 -7550 125 -7530
rect 60 -7560 125 -7550
rect 415 -7530 480 -7520
rect 415 -7550 425 -7530
rect 470 -7550 480 -7530
rect 415 -7560 480 -7550
rect 600 -7530 665 -7520
rect 600 -7550 610 -7530
rect 655 -7550 665 -7530
rect 600 -7560 665 -7550
rect 955 -7530 1020 -7520
rect 955 -7550 965 -7530
rect 1010 -7550 1020 -7530
rect 955 -7560 1020 -7550
rect 1140 -7530 1205 -7520
rect 1140 -7550 1150 -7530
rect 1195 -7550 1205 -7530
rect 1140 -7560 1205 -7550
rect 1495 -7530 1560 -7520
rect 1495 -7550 1505 -7530
rect 1550 -7550 1560 -7530
rect 1495 -7560 1560 -7550
rect 1680 -7530 1745 -7520
rect 1680 -7550 1690 -7530
rect 1735 -7550 1745 -7530
rect 1680 -7560 1745 -7550
rect 2035 -7530 2100 -7520
rect 2035 -7550 2045 -7530
rect 2090 -7550 2100 -7530
rect 2035 -7560 2100 -7550
rect 2220 -7530 2285 -7520
rect 2220 -7550 2230 -7530
rect 2275 -7550 2285 -7530
rect 2220 -7560 2285 -7550
rect 2575 -7530 2640 -7520
rect 2575 -7550 2585 -7530
rect 2630 -7550 2640 -7530
rect 2575 -7560 2640 -7550
rect 2760 -7530 2825 -7520
rect 2760 -7550 2770 -7530
rect 2815 -7550 2825 -7530
rect 2760 -7560 2825 -7550
rect 3115 -7530 3180 -7520
rect 3115 -7550 3125 -7530
rect 3170 -7550 3180 -7530
rect 3115 -7560 3180 -7550
rect 3300 -7530 3365 -7520
rect 3300 -7550 3310 -7530
rect 3355 -7550 3365 -7530
rect 3300 -7560 3365 -7550
rect -40 -7800 0 -7790
rect -40 -7820 -30 -7800
rect -10 -7810 0 -7800
rect 145 -7800 185 -7790
rect 145 -7810 155 -7800
rect -10 -7820 155 -7810
rect 175 -7810 185 -7800
rect 500 -7800 540 -7790
rect 500 -7810 510 -7800
rect 175 -7820 510 -7810
rect 530 -7810 540 -7800
rect 685 -7800 725 -7790
rect 685 -7810 695 -7800
rect 530 -7820 695 -7810
rect 715 -7810 725 -7800
rect 1040 -7800 1080 -7790
rect 1040 -7810 1050 -7800
rect 715 -7820 1050 -7810
rect 1070 -7810 1080 -7800
rect 1225 -7800 1265 -7790
rect 1225 -7810 1235 -7800
rect 1070 -7820 1235 -7810
rect 1255 -7810 1265 -7800
rect 1580 -7800 1620 -7790
rect 1580 -7810 1590 -7800
rect 1255 -7820 1590 -7810
rect 1610 -7810 1620 -7800
rect 1765 -7800 1805 -7790
rect 1765 -7810 1775 -7800
rect 1610 -7820 1775 -7810
rect 1795 -7810 1805 -7800
rect 2120 -7800 2160 -7790
rect 2120 -7810 2130 -7800
rect 1795 -7820 2130 -7810
rect 2150 -7810 2160 -7800
rect 2305 -7800 2345 -7790
rect 2305 -7810 2315 -7800
rect 2150 -7820 2315 -7810
rect 2335 -7810 2345 -7800
rect 2660 -7800 2700 -7790
rect 2660 -7810 2670 -7800
rect 2335 -7820 2670 -7810
rect 2690 -7810 2700 -7800
rect 2845 -7800 2885 -7790
rect 2845 -7810 2855 -7800
rect 2690 -7820 2855 -7810
rect 2875 -7810 2885 -7800
rect 3200 -7800 3240 -7790
rect 3200 -7810 3210 -7800
rect 2875 -7820 3210 -7810
rect 3230 -7810 3240 -7800
rect 3385 -7800 3425 -7790
rect 3385 -7810 3395 -7800
rect 3230 -7820 3395 -7810
rect 3415 -7820 3425 -7800
rect -40 -7830 3425 -7820
rect -125 -8080 -60 -8070
rect -125 -8100 -115 -8080
rect -70 -8090 -60 -8080
rect -20 -8090 0 -7830
rect 60 -8080 125 -8070
rect 60 -8090 70 -8080
rect -70 -8100 70 -8090
rect 115 -8090 125 -8080
rect 415 -8080 480 -8070
rect 415 -8090 425 -8080
rect 115 -8100 425 -8090
rect 470 -8090 480 -8080
rect 600 -8080 665 -8070
rect 600 -8090 610 -8080
rect 470 -8100 610 -8090
rect 655 -8090 665 -8080
rect 955 -8080 1020 -8070
rect 955 -8090 965 -8080
rect 655 -8100 965 -8090
rect 1010 -8090 1020 -8080
rect 1140 -8080 1205 -8070
rect 1140 -8090 1150 -8080
rect 1010 -8100 1150 -8090
rect 1195 -8090 1205 -8080
rect 1495 -8080 1560 -8070
rect 1495 -8090 1505 -8080
rect 1195 -8100 1505 -8090
rect 1550 -8090 1560 -8080
rect 1680 -8080 1745 -8070
rect 1680 -8090 1690 -8080
rect 1550 -8100 1690 -8090
rect 1735 -8090 1745 -8080
rect 2035 -8080 2100 -8070
rect 2035 -8090 2045 -8080
rect 1735 -8100 2045 -8090
rect 2090 -8090 2100 -8080
rect 2220 -8080 2285 -8070
rect 2220 -8090 2230 -8080
rect 2090 -8100 2230 -8090
rect 2275 -8090 2285 -8080
rect 2575 -8080 2640 -8070
rect 2575 -8090 2585 -8080
rect 2275 -8100 2585 -8090
rect 2630 -8090 2640 -8080
rect 2760 -8080 2825 -8070
rect 2760 -8090 2770 -8080
rect 2630 -8100 2770 -8090
rect 2815 -8090 2825 -8080
rect 3115 -8080 3180 -8070
rect 3115 -8090 3125 -8080
rect 2815 -8100 3125 -8090
rect 3170 -8090 3180 -8080
rect 3300 -8080 3365 -8070
rect 3300 -8090 3310 -8080
rect 3170 -8100 3310 -8090
rect 3355 -8100 3365 -8080
rect -125 -8110 3365 -8100
rect 205 -8230 255 -8220
rect 205 -8310 215 -8230
rect 245 -8310 255 -8230
rect 205 -8320 255 -8310
rect 290 -8230 340 -8220
rect 290 -8310 300 -8230
rect 330 -8310 340 -8230
rect 290 -8320 340 -8310
rect 745 -8230 795 -8220
rect 745 -8310 755 -8230
rect 785 -8310 795 -8230
rect 745 -8320 795 -8310
rect 830 -8230 880 -8220
rect 830 -8310 840 -8230
rect 870 -8310 880 -8230
rect 830 -8320 880 -8310
rect 1285 -8230 1335 -8220
rect 1285 -8310 1295 -8230
rect 1325 -8310 1335 -8230
rect 1285 -8320 1335 -8310
rect 1370 -8230 1420 -8220
rect 1370 -8310 1380 -8230
rect 1410 -8310 1420 -8230
rect 1370 -8320 1420 -8310
rect 1825 -8230 1875 -8220
rect 1825 -8310 1835 -8230
rect 1865 -8310 1875 -8230
rect 1825 -8320 1875 -8310
rect 1910 -8230 1960 -8220
rect 1910 -8310 1920 -8230
rect 1950 -8310 1960 -8230
rect 1910 -8320 1960 -8310
rect 2365 -8230 2415 -8220
rect 2365 -8310 2375 -8230
rect 2405 -8310 2415 -8230
rect 2365 -8320 2415 -8310
rect 2450 -8230 2500 -8220
rect 2450 -8310 2460 -8230
rect 2490 -8310 2500 -8230
rect 2450 -8320 2500 -8310
rect 2905 -8230 2955 -8220
rect 2905 -8310 2915 -8230
rect 2945 -8310 2955 -8230
rect 2905 -8320 2955 -8310
rect 2990 -8230 3040 -8220
rect 2990 -8310 3000 -8230
rect 3030 -8310 3040 -8230
rect 2990 -8320 3040 -8310
rect 220 -8340 240 -8320
rect -225 -8360 240 -8340
rect 305 -8380 325 -8320
rect -265 -8400 325 -8380
rect 760 -8420 780 -8320
rect -305 -8440 780 -8420
rect 845 -8460 865 -8320
rect -345 -8480 865 -8460
rect 1300 -8500 1320 -8320
rect -385 -8520 1320 -8500
rect 1385 -8540 1405 -8320
rect -425 -8560 1405 -8540
rect 1840 -8540 1860 -8320
rect 1925 -8500 1945 -8320
rect 2380 -8460 2400 -8320
rect 2465 -8420 2485 -8320
rect 2920 -8380 2940 -8320
rect 3005 -8340 3025 -8320
rect 3800 -8340 3820 3585
rect 3005 -8360 3820 -8340
rect 3840 -8380 3860 3625
rect 2920 -8400 3860 -8380
rect 3880 -8420 3900 3665
rect 2465 -8440 3900 -8420
rect 3920 -8460 3940 3705
rect 2380 -8480 3940 -8460
rect 3960 -8500 3980 3745
rect 1925 -8520 3980 -8500
rect 4000 -8540 4020 3785
rect 1840 -8560 4025 -8540
<< viali >>
rect 215 3460 245 3540
rect 305 3460 335 3540
rect 755 3460 785 3540
rect 845 3460 875 3540
rect 1295 3460 1325 3540
rect 1385 3460 1415 3540
rect 1835 3460 1865 3540
rect 1925 3460 1955 3540
rect 2375 3460 2405 3540
rect 2465 3460 2495 3540
rect 2915 3460 2945 3540
rect 3005 3460 3035 3540
rect -115 2720 -70 2740
rect 70 2720 115 2740
rect 425 2720 470 2740
rect 610 2720 655 2740
rect 965 2720 1010 2740
rect 1150 2720 1195 2740
rect 1505 2720 1550 2740
rect 1690 2720 1735 2740
rect 2045 2720 2090 2740
rect 2230 2720 2275 2740
rect 2585 2720 2630 2740
rect 2770 2720 2815 2740
rect 3125 2720 3170 2740
rect 3310 2720 3355 2740
rect -175 2425 -155 2445
rect 195 2375 250 2405
rect 290 2300 345 2330
rect 735 2375 790 2405
rect 830 2300 885 2330
rect 1275 2375 1330 2405
rect 1370 2300 1425 2330
rect 1815 2375 1870 2405
rect 1910 2300 1965 2330
rect 2355 2375 2410 2405
rect 2450 2300 2505 2330
rect 2895 2375 2950 2405
rect 2990 2300 3045 2330
rect 3750 -2695 3770 -2675
rect -115 -2995 -70 -2975
rect -175 -3290 -155 -3270
rect 290 -7100 345 -7070
rect 195 -7175 250 -7145
rect -175 -7290 -155 -7270
rect 830 -7100 885 -7070
rect 735 -7175 790 -7145
rect 1370 -7100 1425 -7070
rect 1275 -7175 1330 -7145
rect 1910 -7100 1965 -7070
rect 1815 -7175 1870 -7145
rect 2450 -7100 2505 -7070
rect 2355 -7175 2410 -7145
rect 2990 -7100 3045 -7070
rect 2895 -7175 2950 -7145
rect 3435 -7100 3490 -7070
rect -115 -7550 -70 -7530
rect 70 -7550 115 -7530
rect 425 -7550 470 -7530
rect 610 -7550 655 -7530
rect 965 -7550 1010 -7530
rect 1150 -7550 1195 -7530
rect 1505 -7550 1550 -7530
rect 1690 -7550 1735 -7530
rect 2045 -7550 2090 -7530
rect 2230 -7550 2275 -7530
rect 2585 -7550 2630 -7530
rect 2770 -7550 2815 -7530
rect 3125 -7550 3170 -7530
rect 3310 -7550 3355 -7530
rect 215 -8310 245 -8230
rect 300 -8310 330 -8230
rect 755 -8310 785 -8230
rect 840 -8310 870 -8230
rect 1295 -8310 1325 -8230
rect 1380 -8310 1410 -8230
rect 1835 -8310 1865 -8230
rect 1920 -8310 1950 -8230
rect 2375 -8310 2405 -8230
rect 2460 -8310 2490 -8230
rect 2915 -8310 2945 -8230
rect 3000 -8310 3030 -8230
<< metal1 >>
rect 205 3545 255 3550
rect 205 3455 210 3545
rect 250 3455 255 3545
rect 205 3450 255 3455
rect 295 3545 345 3550
rect 295 3455 300 3545
rect 340 3455 345 3545
rect 295 3450 345 3455
rect 745 3545 795 3550
rect 745 3455 750 3545
rect 790 3455 795 3545
rect 745 3450 795 3455
rect 835 3545 885 3550
rect 835 3455 840 3545
rect 880 3455 885 3545
rect 835 3450 885 3455
rect 1285 3545 1335 3550
rect 1285 3455 1290 3545
rect 1330 3455 1335 3545
rect 1285 3450 1335 3455
rect 1375 3545 1425 3550
rect 1375 3455 1380 3545
rect 1420 3455 1425 3545
rect 1375 3450 1425 3455
rect 1825 3545 1875 3550
rect 1825 3455 1830 3545
rect 1870 3455 1875 3545
rect 1825 3450 1875 3455
rect 1915 3545 1965 3550
rect 1915 3455 1920 3545
rect 1960 3455 1965 3545
rect 1915 3450 1965 3455
rect 2365 3545 2415 3550
rect 2365 3455 2370 3545
rect 2410 3455 2415 3545
rect 2365 3450 2415 3455
rect 2455 3545 2505 3550
rect 2455 3455 2460 3545
rect 2500 3455 2505 3545
rect 2455 3450 2505 3455
rect 2905 3545 2955 3550
rect 2905 3455 2910 3545
rect 2950 3455 2955 3545
rect 2905 3450 2955 3455
rect 2995 3545 3045 3550
rect 2995 3455 3000 3545
rect 3040 3455 3045 3545
rect 2995 3450 3045 3455
rect -180 3320 4060 3340
rect -180 2750 -160 3320
rect -130 2750 -55 2755
rect -180 2740 -55 2750
rect -180 2720 -115 2740
rect -70 2720 -55 2740
rect -180 2710 -55 2720
rect -130 2705 -55 2710
rect 55 2740 130 2755
rect 55 2720 70 2740
rect 115 2720 130 2740
rect 55 2705 130 2720
rect 360 2750 380 3320
rect 410 2750 485 2755
rect 360 2740 485 2750
rect 360 2720 425 2740
rect 470 2720 485 2740
rect 360 2710 485 2720
rect 410 2705 485 2710
rect 595 2740 670 2755
rect 595 2720 610 2740
rect 655 2720 670 2740
rect 595 2705 670 2720
rect 900 2750 920 3320
rect 950 2750 1025 2755
rect 900 2740 1025 2750
rect 900 2720 965 2740
rect 1010 2720 1025 2740
rect 900 2710 1025 2720
rect 950 2705 1025 2710
rect 1135 2740 1210 2755
rect 1135 2720 1150 2740
rect 1195 2720 1210 2740
rect 1135 2705 1210 2720
rect 1440 2750 1460 3320
rect 1490 2750 1565 2755
rect 1440 2740 1565 2750
rect 1440 2720 1505 2740
rect 1550 2720 1565 2740
rect 1440 2710 1565 2720
rect 1490 2705 1565 2710
rect 1675 2740 1750 2755
rect 1675 2720 1690 2740
rect 1735 2720 1750 2740
rect 1675 2705 1750 2720
rect 1980 2750 2000 3320
rect 2030 2750 2105 2755
rect 1980 2740 2105 2750
rect 1980 2720 2045 2740
rect 2090 2720 2105 2740
rect 1980 2710 2105 2720
rect 2030 2705 2105 2710
rect 2215 2740 2290 2755
rect 2215 2720 2230 2740
rect 2275 2720 2290 2740
rect 2215 2705 2290 2720
rect 2520 2750 2540 3320
rect 2570 2750 2645 2755
rect 2520 2740 2645 2750
rect 2520 2720 2585 2740
rect 2630 2720 2645 2740
rect 2520 2710 2645 2720
rect 2570 2705 2645 2710
rect 2755 2740 2830 2755
rect 2755 2720 2770 2740
rect 2815 2720 2830 2740
rect 2755 2705 2830 2720
rect 3060 2750 3080 3320
rect 3110 2750 3185 2755
rect 3060 2740 3185 2750
rect 3060 2720 3125 2740
rect 3170 2720 3185 2740
rect 3060 2710 3185 2720
rect 3110 2705 3185 2710
rect 3295 2740 3370 2755
rect 3295 2720 3310 2740
rect 3355 2720 3370 2740
rect 3295 2705 3370 2720
rect -205 2445 -145 2455
rect -205 2425 -175 2445
rect -155 2425 -145 2445
rect -205 2415 -145 2425
rect -205 -2975 -185 2415
rect 185 2410 260 2415
rect 185 2370 190 2410
rect 255 2370 260 2410
rect 185 2365 260 2370
rect 725 2410 800 2415
rect 725 2370 730 2410
rect 795 2370 800 2410
rect 725 2365 800 2370
rect 1265 2410 1340 2415
rect 1265 2370 1270 2410
rect 1335 2370 1340 2410
rect 1265 2365 1340 2370
rect 1805 2410 1880 2415
rect 1805 2370 1810 2410
rect 1875 2370 1880 2410
rect 1805 2365 1880 2370
rect 2345 2410 2420 2415
rect 2345 2370 2350 2410
rect 2415 2370 2420 2410
rect 2345 2365 2420 2370
rect 2885 2410 2960 2415
rect 2885 2370 2890 2410
rect 2955 2370 2960 2410
rect 2885 2365 2960 2370
rect 280 2335 355 2340
rect 280 2295 285 2335
rect 350 2295 355 2335
rect 280 2290 355 2295
rect 820 2335 895 2340
rect 820 2295 825 2335
rect 890 2295 895 2335
rect 820 2290 895 2295
rect 1360 2335 1435 2340
rect 1360 2295 1365 2335
rect 1430 2295 1435 2335
rect 1360 2290 1435 2295
rect 1900 2335 1975 2340
rect 1900 2295 1905 2335
rect 1970 2295 1975 2335
rect 1900 2290 1975 2295
rect 2440 2335 2515 2340
rect 2440 2295 2445 2335
rect 2510 2295 2515 2335
rect 2440 2290 2515 2295
rect 2980 2335 3055 2340
rect 2980 2295 2985 2335
rect 3050 2295 3055 2335
rect 2980 2290 3055 2295
rect 3740 -2670 3780 -2665
rect 3740 -2700 3745 -2670
rect 3775 -2700 3780 -2670
rect 3740 -2705 3780 -2700
rect -130 -2975 -55 -2960
rect -450 -2995 -115 -2975
rect -70 -2995 -55 -2975
rect -205 -3260 -185 -2995
rect -130 -3010 -55 -2995
rect -205 -3270 -145 -3260
rect -450 -3290 -175 -3270
rect -155 -3290 -145 -3270
rect -205 -3300 -145 -3290
rect -205 -7260 -185 -3300
rect 280 -7065 355 -7060
rect 280 -7105 285 -7065
rect 350 -7105 355 -7065
rect 280 -7110 355 -7105
rect 820 -7065 895 -7060
rect 820 -7105 825 -7065
rect 890 -7105 895 -7065
rect 820 -7110 895 -7105
rect 1360 -7065 1435 -7060
rect 1360 -7105 1365 -7065
rect 1430 -7105 1435 -7065
rect 1360 -7110 1435 -7105
rect 1900 -7065 1975 -7060
rect 1900 -7105 1905 -7065
rect 1970 -7105 1975 -7065
rect 1900 -7110 1975 -7105
rect 2440 -7065 2515 -7060
rect 2440 -7105 2445 -7065
rect 2510 -7105 2515 -7065
rect 2440 -7110 2515 -7105
rect 2980 -7065 3055 -7060
rect 2980 -7105 2985 -7065
rect 3050 -7105 3055 -7065
rect 2980 -7110 3055 -7105
rect 3425 -7065 3500 -7060
rect 3425 -7105 3430 -7065
rect 3495 -7105 3500 -7065
rect 3425 -7110 3500 -7105
rect 185 -7140 260 -7135
rect 185 -7180 190 -7140
rect 255 -7180 260 -7140
rect 185 -7185 260 -7180
rect 725 -7140 800 -7135
rect 725 -7180 730 -7140
rect 795 -7180 800 -7140
rect 725 -7185 800 -7180
rect 1265 -7140 1340 -7135
rect 1265 -7180 1270 -7140
rect 1335 -7180 1340 -7140
rect 1265 -7185 1340 -7180
rect 1805 -7140 1880 -7135
rect 1805 -7180 1810 -7140
rect 1875 -7180 1880 -7140
rect 1805 -7185 1880 -7180
rect 2345 -7140 2420 -7135
rect 2345 -7180 2350 -7140
rect 2415 -7180 2420 -7140
rect 2345 -7185 2420 -7180
rect 2885 -7140 2960 -7135
rect 2885 -7180 2890 -7140
rect 2955 -7180 2960 -7140
rect 2885 -7185 2960 -7180
rect -205 -7270 -145 -7260
rect -440 -7290 -175 -7270
rect -155 -7290 -145 -7270
rect -185 -7300 -145 -7290
rect 55 -7520 130 -7515
rect 410 -7520 485 -7515
rect 950 -7520 1025 -7515
rect 1490 -7520 1565 -7515
rect 2030 -7520 2105 -7515
rect 2570 -7520 2645 -7515
rect 3110 -7520 3185 -7515
rect -185 -7530 -55 -7520
rect -185 -7550 -115 -7530
rect -70 -7550 -55 -7530
rect -185 -7560 -55 -7550
rect 55 -7560 60 -7520
rect 125 -7560 130 -7520
rect -185 -8130 -165 -7560
rect 55 -7565 130 -7560
rect 355 -7530 485 -7520
rect 355 -7550 425 -7530
rect 470 -7550 485 -7530
rect 355 -7560 485 -7550
rect 595 -7560 600 -7520
rect 665 -7560 670 -7520
rect 895 -7530 1025 -7520
rect 895 -7550 965 -7530
rect 1010 -7550 1025 -7530
rect 895 -7560 1025 -7550
rect 1135 -7560 1140 -7520
rect 1205 -7560 1210 -7520
rect 1435 -7530 1565 -7520
rect 1435 -7550 1505 -7530
rect 1550 -7550 1565 -7530
rect 1435 -7560 1565 -7550
rect 1675 -7560 1680 -7520
rect 1745 -7560 1750 -7520
rect 1975 -7530 2105 -7520
rect 1975 -7550 2045 -7530
rect 2090 -7550 2105 -7530
rect 1975 -7560 2105 -7550
rect 2215 -7560 2220 -7520
rect 2285 -7560 2290 -7520
rect 2515 -7530 2645 -7520
rect 2515 -7550 2585 -7530
rect 2630 -7550 2645 -7530
rect 2515 -7560 2645 -7550
rect 2755 -7560 2760 -7520
rect 2825 -7560 2830 -7520
rect 3055 -7530 3185 -7520
rect 3055 -7550 3125 -7530
rect 3170 -7550 3185 -7530
rect 3055 -7560 3185 -7550
rect 3295 -7560 3300 -7520
rect 3365 -7560 3370 -7520
rect 355 -8130 375 -7560
rect 410 -7565 485 -7560
rect 895 -8130 915 -7560
rect 950 -7565 1025 -7560
rect 1435 -8130 1455 -7560
rect 1490 -7565 1565 -7560
rect 1975 -8130 1995 -7560
rect 2030 -7565 2105 -7560
rect 2515 -8130 2535 -7560
rect 2570 -7565 2645 -7560
rect 3055 -8130 3075 -7560
rect 3110 -7565 3185 -7560
rect 4040 -8130 4060 3320
rect -185 -8150 4340 -8130
rect 205 -8225 255 -8220
rect 205 -8315 210 -8225
rect 250 -8315 255 -8225
rect 205 -8320 255 -8315
rect 290 -8225 340 -8220
rect 290 -8315 295 -8225
rect 335 -8315 340 -8225
rect 290 -8320 340 -8315
rect 745 -8225 795 -8220
rect 745 -8315 750 -8225
rect 790 -8315 795 -8225
rect 745 -8320 795 -8315
rect 830 -8225 880 -8220
rect 830 -8315 835 -8225
rect 875 -8315 880 -8225
rect 830 -8320 880 -8315
rect 1285 -8225 1335 -8220
rect 1285 -8315 1290 -8225
rect 1330 -8315 1335 -8225
rect 1285 -8320 1335 -8315
rect 1370 -8225 1420 -8220
rect 1370 -8315 1375 -8225
rect 1415 -8315 1420 -8225
rect 1370 -8320 1420 -8315
rect 1825 -8225 1875 -8220
rect 1825 -8315 1830 -8225
rect 1870 -8315 1875 -8225
rect 1825 -8320 1875 -8315
rect 1910 -8225 1960 -8220
rect 1910 -8315 1915 -8225
rect 1955 -8315 1960 -8225
rect 1910 -8320 1960 -8315
rect 2365 -8225 2415 -8220
rect 2365 -8315 2370 -8225
rect 2410 -8315 2415 -8225
rect 2365 -8320 2415 -8315
rect 2450 -8225 2500 -8220
rect 2450 -8315 2455 -8225
rect 2495 -8315 2500 -8225
rect 2450 -8320 2500 -8315
rect 2905 -8225 2955 -8220
rect 2905 -8315 2910 -8225
rect 2950 -8315 2955 -8225
rect 2905 -8320 2955 -8315
rect 2990 -8225 3040 -8220
rect 2990 -8315 2995 -8225
rect 3035 -8315 3040 -8225
rect 2990 -8320 3040 -8315
<< via1 >>
rect 210 3540 250 3545
rect 210 3460 215 3540
rect 215 3460 245 3540
rect 245 3460 250 3540
rect 210 3455 250 3460
rect 300 3540 340 3545
rect 300 3460 305 3540
rect 305 3460 335 3540
rect 335 3460 340 3540
rect 300 3455 340 3460
rect 750 3540 790 3545
rect 750 3460 755 3540
rect 755 3460 785 3540
rect 785 3460 790 3540
rect 750 3455 790 3460
rect 840 3540 880 3545
rect 840 3460 845 3540
rect 845 3460 875 3540
rect 875 3460 880 3540
rect 840 3455 880 3460
rect 1290 3540 1330 3545
rect 1290 3460 1295 3540
rect 1295 3460 1325 3540
rect 1325 3460 1330 3540
rect 1290 3455 1330 3460
rect 1380 3540 1420 3545
rect 1380 3460 1385 3540
rect 1385 3460 1415 3540
rect 1415 3460 1420 3540
rect 1380 3455 1420 3460
rect 1830 3540 1870 3545
rect 1830 3460 1835 3540
rect 1835 3460 1865 3540
rect 1865 3460 1870 3540
rect 1830 3455 1870 3460
rect 1920 3540 1960 3545
rect 1920 3460 1925 3540
rect 1925 3460 1955 3540
rect 1955 3460 1960 3540
rect 1920 3455 1960 3460
rect 2370 3540 2410 3545
rect 2370 3460 2375 3540
rect 2375 3460 2405 3540
rect 2405 3460 2410 3540
rect 2370 3455 2410 3460
rect 2460 3540 2500 3545
rect 2460 3460 2465 3540
rect 2465 3460 2495 3540
rect 2495 3460 2500 3540
rect 2460 3455 2500 3460
rect 2910 3540 2950 3545
rect 2910 3460 2915 3540
rect 2915 3460 2945 3540
rect 2945 3460 2950 3540
rect 2910 3455 2950 3460
rect 3000 3540 3040 3545
rect 3000 3460 3005 3540
rect 3005 3460 3035 3540
rect 3035 3460 3040 3540
rect 3000 3455 3040 3460
rect 190 2405 255 2410
rect 190 2375 195 2405
rect 195 2375 250 2405
rect 250 2375 255 2405
rect 190 2370 255 2375
rect 730 2405 795 2410
rect 730 2375 735 2405
rect 735 2375 790 2405
rect 790 2375 795 2405
rect 730 2370 795 2375
rect 1270 2405 1335 2410
rect 1270 2375 1275 2405
rect 1275 2375 1330 2405
rect 1330 2375 1335 2405
rect 1270 2370 1335 2375
rect 1810 2405 1875 2410
rect 1810 2375 1815 2405
rect 1815 2375 1870 2405
rect 1870 2375 1875 2405
rect 1810 2370 1875 2375
rect 2350 2405 2415 2410
rect 2350 2375 2355 2405
rect 2355 2375 2410 2405
rect 2410 2375 2415 2405
rect 2350 2370 2415 2375
rect 2890 2405 2955 2410
rect 2890 2375 2895 2405
rect 2895 2375 2950 2405
rect 2950 2375 2955 2405
rect 2890 2370 2955 2375
rect 285 2330 350 2335
rect 285 2300 290 2330
rect 290 2300 345 2330
rect 345 2300 350 2330
rect 285 2295 350 2300
rect 825 2330 890 2335
rect 825 2300 830 2330
rect 830 2300 885 2330
rect 885 2300 890 2330
rect 825 2295 890 2300
rect 1365 2330 1430 2335
rect 1365 2300 1370 2330
rect 1370 2300 1425 2330
rect 1425 2300 1430 2330
rect 1365 2295 1430 2300
rect 1905 2330 1970 2335
rect 1905 2300 1910 2330
rect 1910 2300 1965 2330
rect 1965 2300 1970 2330
rect 1905 2295 1970 2300
rect 2445 2330 2510 2335
rect 2445 2300 2450 2330
rect 2450 2300 2505 2330
rect 2505 2300 2510 2330
rect 2445 2295 2510 2300
rect 2985 2330 3050 2335
rect 2985 2300 2990 2330
rect 2990 2300 3045 2330
rect 3045 2300 3050 2330
rect 2985 2295 3050 2300
rect 3745 -2675 3775 -2670
rect 3745 -2695 3750 -2675
rect 3750 -2695 3770 -2675
rect 3770 -2695 3775 -2675
rect 3745 -2700 3775 -2695
rect 285 -7070 350 -7065
rect 285 -7100 290 -7070
rect 290 -7100 345 -7070
rect 345 -7100 350 -7070
rect 285 -7105 350 -7100
rect 825 -7070 890 -7065
rect 825 -7100 830 -7070
rect 830 -7100 885 -7070
rect 885 -7100 890 -7070
rect 825 -7105 890 -7100
rect 1365 -7070 1430 -7065
rect 1365 -7100 1370 -7070
rect 1370 -7100 1425 -7070
rect 1425 -7100 1430 -7070
rect 1365 -7105 1430 -7100
rect 1905 -7070 1970 -7065
rect 1905 -7100 1910 -7070
rect 1910 -7100 1965 -7070
rect 1965 -7100 1970 -7070
rect 1905 -7105 1970 -7100
rect 2445 -7070 2510 -7065
rect 2445 -7100 2450 -7070
rect 2450 -7100 2505 -7070
rect 2505 -7100 2510 -7070
rect 2445 -7105 2510 -7100
rect 2985 -7070 3050 -7065
rect 2985 -7100 2990 -7070
rect 2990 -7100 3045 -7070
rect 3045 -7100 3050 -7070
rect 2985 -7105 3050 -7100
rect 3430 -7070 3495 -7065
rect 3430 -7100 3435 -7070
rect 3435 -7100 3490 -7070
rect 3490 -7100 3495 -7070
rect 3430 -7105 3495 -7100
rect 190 -7145 255 -7140
rect 190 -7175 195 -7145
rect 195 -7175 250 -7145
rect 250 -7175 255 -7145
rect 190 -7180 255 -7175
rect 730 -7145 795 -7140
rect 730 -7175 735 -7145
rect 735 -7175 790 -7145
rect 790 -7175 795 -7145
rect 730 -7180 795 -7175
rect 1270 -7145 1335 -7140
rect 1270 -7175 1275 -7145
rect 1275 -7175 1330 -7145
rect 1330 -7175 1335 -7145
rect 1270 -7180 1335 -7175
rect 1810 -7145 1875 -7140
rect 1810 -7175 1815 -7145
rect 1815 -7175 1870 -7145
rect 1870 -7175 1875 -7145
rect 1810 -7180 1875 -7175
rect 2350 -7145 2415 -7140
rect 2350 -7175 2355 -7145
rect 2355 -7175 2410 -7145
rect 2410 -7175 2415 -7145
rect 2350 -7180 2415 -7175
rect 2890 -7145 2955 -7140
rect 2890 -7175 2895 -7145
rect 2895 -7175 2950 -7145
rect 2950 -7175 2955 -7145
rect 2890 -7180 2955 -7175
rect 60 -7530 125 -7520
rect 60 -7550 70 -7530
rect 70 -7550 115 -7530
rect 115 -7550 125 -7530
rect 60 -7560 125 -7550
rect 600 -7530 665 -7520
rect 600 -7550 610 -7530
rect 610 -7550 655 -7530
rect 655 -7550 665 -7530
rect 600 -7560 665 -7550
rect 1140 -7530 1205 -7520
rect 1140 -7550 1150 -7530
rect 1150 -7550 1195 -7530
rect 1195 -7550 1205 -7530
rect 1140 -7560 1205 -7550
rect 1680 -7530 1745 -7520
rect 1680 -7550 1690 -7530
rect 1690 -7550 1735 -7530
rect 1735 -7550 1745 -7530
rect 1680 -7560 1745 -7550
rect 2220 -7530 2285 -7520
rect 2220 -7550 2230 -7530
rect 2230 -7550 2275 -7530
rect 2275 -7550 2285 -7530
rect 2220 -7560 2285 -7550
rect 2760 -7530 2825 -7520
rect 2760 -7550 2770 -7530
rect 2770 -7550 2815 -7530
rect 2815 -7550 2825 -7530
rect 2760 -7560 2825 -7550
rect 3300 -7530 3365 -7520
rect 3300 -7550 3310 -7530
rect 3310 -7550 3355 -7530
rect 3355 -7550 3365 -7530
rect 3300 -7560 3365 -7550
rect 210 -8230 250 -8225
rect 210 -8310 215 -8230
rect 215 -8310 245 -8230
rect 245 -8310 250 -8230
rect 210 -8315 250 -8310
rect 295 -8230 335 -8225
rect 295 -8310 300 -8230
rect 300 -8310 330 -8230
rect 330 -8310 335 -8230
rect 295 -8315 335 -8310
rect 750 -8230 790 -8225
rect 750 -8310 755 -8230
rect 755 -8310 785 -8230
rect 785 -8310 790 -8230
rect 750 -8315 790 -8310
rect 835 -8230 875 -8225
rect 835 -8310 840 -8230
rect 840 -8310 870 -8230
rect 870 -8310 875 -8230
rect 835 -8315 875 -8310
rect 1290 -8230 1330 -8225
rect 1290 -8310 1295 -8230
rect 1295 -8310 1325 -8230
rect 1325 -8310 1330 -8230
rect 1290 -8315 1330 -8310
rect 1375 -8230 1415 -8225
rect 1375 -8310 1380 -8230
rect 1380 -8310 1410 -8230
rect 1410 -8310 1415 -8230
rect 1375 -8315 1415 -8310
rect 1830 -8230 1870 -8225
rect 1830 -8310 1835 -8230
rect 1835 -8310 1865 -8230
rect 1865 -8310 1870 -8230
rect 1830 -8315 1870 -8310
rect 1915 -8230 1955 -8225
rect 1915 -8310 1920 -8230
rect 1920 -8310 1950 -8230
rect 1950 -8310 1955 -8230
rect 1915 -8315 1955 -8310
rect 2370 -8230 2410 -8225
rect 2370 -8310 2375 -8230
rect 2375 -8310 2405 -8230
rect 2405 -8310 2410 -8230
rect 2370 -8315 2410 -8310
rect 2455 -8230 2495 -8225
rect 2455 -8310 2460 -8230
rect 2460 -8310 2490 -8230
rect 2490 -8310 2495 -8230
rect 2455 -8315 2495 -8310
rect 2910 -8230 2950 -8225
rect 2910 -8310 2915 -8230
rect 2915 -8310 2945 -8230
rect 2945 -8310 2950 -8230
rect 2910 -8315 2950 -8310
rect 2995 -8230 3035 -8225
rect 2995 -8310 3000 -8230
rect 3000 -8310 3030 -8230
rect 3030 -8310 3035 -8230
rect 2995 -8315 3035 -8310
<< metal2 >>
rect 205 3545 255 3550
rect 205 3455 210 3545
rect 250 3455 255 3545
rect 205 3450 255 3455
rect 295 3545 345 3550
rect 295 3455 300 3545
rect 340 3455 345 3545
rect 295 3450 345 3455
rect 745 3545 795 3550
rect 745 3455 750 3545
rect 790 3455 795 3545
rect 745 3450 795 3455
rect 835 3545 885 3550
rect 835 3455 840 3545
rect 880 3455 885 3545
rect 835 3450 885 3455
rect 1285 3545 1335 3550
rect 1285 3455 1290 3545
rect 1330 3455 1335 3545
rect 1285 3450 1335 3455
rect 1375 3545 1425 3550
rect 1375 3455 1380 3545
rect 1420 3455 1425 3545
rect 1375 3450 1425 3455
rect 1825 3545 1875 3550
rect 1825 3455 1830 3545
rect 1870 3455 1875 3545
rect 1825 3450 1875 3455
rect 1915 3545 1965 3550
rect 1915 3455 1920 3545
rect 1960 3455 1965 3545
rect 1915 3450 1965 3455
rect 2365 3545 2415 3550
rect 2365 3455 2370 3545
rect 2410 3455 2415 3545
rect 2365 3450 2415 3455
rect 2455 3545 2505 3550
rect 2455 3455 2460 3545
rect 2500 3455 2505 3545
rect 2455 3450 2505 3455
rect 2905 3545 2955 3550
rect 2905 3455 2910 3545
rect 2950 3455 2955 3545
rect 2905 3450 2955 3455
rect 2995 3545 3045 3550
rect 2995 3455 3000 3545
rect 3040 3455 3045 3545
rect 2995 3450 3045 3455
rect 10 3360 4100 3380
rect 10 2745 30 3360
rect 55 2745 130 2755
rect 10 2715 130 2745
rect 550 2745 570 3360
rect 595 2745 670 2755
rect 550 2715 670 2745
rect 1090 2745 1110 3360
rect 1135 2745 1210 2755
rect 1090 2715 1210 2745
rect 1630 2745 1650 3360
rect 1675 2745 1750 2755
rect 1630 2715 1750 2745
rect 2170 2745 2190 3360
rect 2215 2745 2290 2755
rect 2170 2715 2290 2745
rect 2710 2745 2730 3360
rect 2755 2745 2830 2755
rect 2710 2715 2830 2745
rect 3250 2745 3270 3360
rect 3295 2745 3370 2755
rect 3250 2715 3370 2745
rect 55 2705 130 2715
rect 595 2705 670 2715
rect 1135 2705 1210 2715
rect 1675 2705 1750 2715
rect 2215 2705 2290 2715
rect 2755 2705 2830 2715
rect 3295 2705 3370 2715
rect 185 2410 260 2415
rect 185 2370 190 2410
rect 255 2370 260 2410
rect 185 2365 260 2370
rect 725 2410 800 2415
rect 725 2370 730 2410
rect 795 2370 800 2410
rect 725 2365 800 2370
rect 1265 2410 1340 2415
rect 1265 2370 1270 2410
rect 1335 2370 1340 2410
rect 1265 2365 1340 2370
rect 1805 2410 1880 2415
rect 1805 2370 1810 2410
rect 1875 2370 1880 2410
rect 1805 2365 1880 2370
rect 2345 2410 2420 2415
rect 2345 2370 2350 2410
rect 2415 2370 2420 2410
rect 2345 2365 2420 2370
rect 2885 2410 2960 2415
rect 2885 2370 2890 2410
rect 2955 2370 2960 2410
rect 2885 2365 2960 2370
rect 280 2335 355 2340
rect 280 2295 285 2335
rect 350 2295 355 2335
rect 280 2290 355 2295
rect 820 2335 895 2340
rect 820 2295 825 2335
rect 890 2295 895 2335
rect 820 2290 895 2295
rect 1360 2335 1435 2340
rect 1360 2295 1365 2335
rect 1430 2295 1435 2335
rect 1360 2290 1435 2295
rect 1900 2335 1975 2340
rect 1900 2295 1905 2335
rect 1970 2295 1975 2335
rect 1900 2290 1975 2295
rect 2440 2335 2515 2340
rect 2440 2295 2445 2335
rect 2510 2295 2515 2335
rect 2440 2290 2515 2295
rect 2980 2335 3055 2340
rect 2980 2295 2985 2335
rect 3050 2295 3055 2335
rect 2980 2290 3055 2295
rect -450 -2650 3760 -2625
rect 3740 -2665 3760 -2650
rect 3740 -2670 3780 -2665
rect 3740 -2700 3745 -2670
rect 3775 -2700 3780 -2670
rect 3740 -2705 3780 -2700
rect 280 -7065 355 -7060
rect 280 -7105 285 -7065
rect 350 -7105 355 -7065
rect 280 -7110 355 -7105
rect 820 -7065 895 -7060
rect 820 -7105 825 -7065
rect 890 -7105 895 -7065
rect 820 -7110 895 -7105
rect 1360 -7065 1435 -7060
rect 1360 -7105 1365 -7065
rect 1430 -7105 1435 -7065
rect 1360 -7110 1435 -7105
rect 1900 -7065 1975 -7060
rect 1900 -7105 1905 -7065
rect 1970 -7105 1975 -7065
rect 1900 -7110 1975 -7105
rect 2440 -7065 2515 -7060
rect 2440 -7105 2445 -7065
rect 2510 -7105 2515 -7065
rect 2440 -7110 2515 -7105
rect 2980 -7065 3055 -7060
rect 2980 -7105 2985 -7065
rect 3050 -7105 3055 -7065
rect 2980 -7110 3055 -7105
rect 3425 -7065 3500 -7060
rect 3425 -7105 3430 -7065
rect 3495 -7105 3500 -7065
rect 3425 -7110 3500 -7105
rect 185 -7140 260 -7135
rect 185 -7180 190 -7140
rect 255 -7180 260 -7140
rect 185 -7185 260 -7180
rect 725 -7140 800 -7135
rect 725 -7180 730 -7140
rect 795 -7180 800 -7140
rect 725 -7185 800 -7180
rect 1265 -7140 1340 -7135
rect 1265 -7180 1270 -7140
rect 1335 -7180 1340 -7140
rect 1265 -7185 1340 -7180
rect 1805 -7140 1880 -7135
rect 1805 -7180 1810 -7140
rect 1875 -7180 1880 -7140
rect 1805 -7185 1880 -7180
rect 2345 -7140 2420 -7135
rect 2345 -7180 2350 -7140
rect 2415 -7180 2420 -7140
rect 2345 -7185 2420 -7180
rect 2885 -7140 2960 -7135
rect 2885 -7180 2890 -7140
rect 2955 -7180 2960 -7140
rect 2885 -7185 2960 -7180
rect 55 -7520 130 -7515
rect 595 -7520 670 -7515
rect 1135 -7520 1210 -7515
rect 1675 -7520 1750 -7515
rect 2215 -7520 2290 -7515
rect 2755 -7520 2830 -7515
rect 3295 -7520 3370 -7515
rect 5 -7560 60 -7520
rect 125 -7560 130 -7520
rect 5 -8170 25 -7560
rect 55 -7565 130 -7560
rect 550 -7560 600 -7520
rect 665 -7560 670 -7520
rect 550 -8170 570 -7560
rect 595 -7565 670 -7560
rect 1090 -7560 1140 -7520
rect 1205 -7560 1210 -7520
rect 1090 -8170 1110 -7560
rect 1135 -7565 1210 -7560
rect 1630 -7560 1680 -7520
rect 1745 -7560 1750 -7520
rect 1630 -8170 1650 -7560
rect 1675 -7565 1750 -7560
rect 2170 -7560 2220 -7520
rect 2285 -7560 2290 -7520
rect 2170 -8170 2190 -7560
rect 2215 -7565 2290 -7560
rect 2710 -7560 2760 -7520
rect 2825 -7560 2830 -7520
rect 2710 -8170 2730 -7560
rect 2755 -7565 2830 -7560
rect 3250 -7560 3300 -7520
rect 3365 -7560 3370 -7520
rect 3250 -8170 3270 -7560
rect 3295 -7565 3370 -7560
rect 4080 -8170 4100 3360
rect 5 -8195 4340 -8170
rect 205 -8225 255 -8220
rect 205 -8315 210 -8225
rect 250 -8315 255 -8225
rect 205 -8320 255 -8315
rect 290 -8225 340 -8220
rect 290 -8315 295 -8225
rect 335 -8315 340 -8225
rect 290 -8320 340 -8315
rect 745 -8225 795 -8220
rect 745 -8315 750 -8225
rect 790 -8315 795 -8225
rect 745 -8320 795 -8315
rect 830 -8225 880 -8220
rect 830 -8315 835 -8225
rect 875 -8315 880 -8225
rect 830 -8320 880 -8315
rect 1285 -8225 1335 -8220
rect 1285 -8315 1290 -8225
rect 1330 -8315 1335 -8225
rect 1285 -8320 1335 -8315
rect 1370 -8225 1420 -8220
rect 1370 -8315 1375 -8225
rect 1415 -8315 1420 -8225
rect 1370 -8320 1420 -8315
rect 1825 -8225 1875 -8220
rect 1825 -8315 1830 -8225
rect 1870 -8315 1875 -8225
rect 1825 -8320 1875 -8315
rect 1910 -8225 1960 -8220
rect 1910 -8315 1915 -8225
rect 1955 -8315 1960 -8225
rect 1910 -8320 1960 -8315
rect 2365 -8225 2415 -8220
rect 2365 -8315 2370 -8225
rect 2410 -8315 2415 -8225
rect 2365 -8320 2415 -8315
rect 2450 -8225 2500 -8220
rect 2450 -8315 2455 -8225
rect 2495 -8315 2500 -8225
rect 2450 -8320 2500 -8315
rect 2905 -8225 2955 -8220
rect 2905 -8315 2910 -8225
rect 2950 -8315 2955 -8225
rect 2905 -8320 2955 -8315
rect 2990 -8225 3040 -8220
rect 2990 -8315 2995 -8225
rect 3035 -8315 3040 -8225
rect 2990 -8320 3040 -8315
<< via2 >>
rect 210 3455 250 3545
rect 300 3455 340 3545
rect 750 3455 790 3545
rect 840 3455 880 3545
rect 1290 3455 1330 3545
rect 1380 3455 1420 3545
rect 1830 3455 1870 3545
rect 1920 3455 1960 3545
rect 2370 3455 2410 3545
rect 2460 3455 2500 3545
rect 2910 3455 2950 3545
rect 3000 3455 3040 3545
rect 190 2370 255 2410
rect 730 2370 795 2410
rect 1270 2370 1335 2410
rect 1810 2370 1875 2410
rect 2350 2370 2415 2410
rect 2890 2370 2955 2410
rect 285 2295 350 2335
rect 825 2295 890 2335
rect 1365 2295 1430 2335
rect 1905 2295 1970 2335
rect 2445 2295 2510 2335
rect 2985 2295 3050 2335
rect 285 -7105 350 -7065
rect 825 -7105 890 -7065
rect 1365 -7105 1430 -7065
rect 1905 -7105 1970 -7065
rect 2445 -7105 2510 -7065
rect 2985 -7105 3050 -7065
rect 3430 -7105 3495 -7065
rect 190 -7180 255 -7140
rect 730 -7180 795 -7140
rect 1270 -7180 1335 -7140
rect 1810 -7180 1875 -7140
rect 2350 -7180 2415 -7140
rect 2890 -7180 2955 -7140
rect 210 -8315 250 -8225
rect 295 -8315 335 -8225
rect 750 -8315 790 -8225
rect 835 -8315 875 -8225
rect 1290 -8315 1330 -8225
rect 1375 -8315 1415 -8225
rect 1830 -8315 1870 -8225
rect 1915 -8315 1955 -8225
rect 2370 -8315 2410 -8225
rect 2455 -8315 2495 -8225
rect 2910 -8315 2950 -8225
rect 2995 -8315 3035 -8225
<< metal3 >>
rect 205 3545 255 3550
rect 205 3455 210 3545
rect 250 3455 255 3545
rect 205 3450 255 3455
rect 295 3545 345 3550
rect 295 3455 300 3545
rect 340 3455 345 3545
rect 295 3450 345 3455
rect 745 3545 795 3550
rect 745 3455 750 3545
rect 790 3455 795 3545
rect 745 3450 795 3455
rect 835 3545 885 3550
rect 835 3455 840 3545
rect 880 3455 885 3545
rect 835 3450 885 3455
rect 1285 3545 1335 3550
rect 1285 3455 1290 3545
rect 1330 3455 1335 3545
rect 1285 3450 1335 3455
rect 1375 3545 1425 3550
rect 1375 3455 1380 3545
rect 1420 3455 1425 3545
rect 1375 3450 1425 3455
rect 1825 3545 1875 3550
rect 1825 3455 1830 3545
rect 1870 3455 1875 3545
rect 1825 3450 1875 3455
rect 1915 3545 1965 3550
rect 1915 3455 1920 3545
rect 1960 3455 1965 3545
rect 1915 3450 1965 3455
rect 2365 3545 2415 3550
rect 2365 3455 2370 3545
rect 2410 3455 2415 3545
rect 2365 3450 2415 3455
rect 2455 3545 2505 3550
rect 2455 3455 2460 3545
rect 2500 3455 2505 3545
rect 2455 3450 2505 3455
rect 2905 3545 2955 3550
rect 2905 3455 2910 3545
rect 2950 3455 2955 3545
rect 2905 3450 2955 3455
rect 2995 3545 3045 3550
rect 2995 3455 3000 3545
rect 3040 3455 3045 3545
rect 2995 3450 3045 3455
rect 215 3060 245 3450
rect 215 2415 245 3030
rect 185 2410 260 2415
rect 185 2370 190 2410
rect 255 2370 260 2410
rect 185 2365 260 2370
rect 305 2340 335 3450
rect 755 3060 785 3450
rect 755 2415 785 3030
rect 725 2410 800 2415
rect 725 2370 730 2410
rect 795 2370 800 2410
rect 725 2365 800 2370
rect 845 2340 875 3450
rect 1295 3060 1325 3450
rect 1295 2415 1325 3030
rect 1265 2410 1340 2415
rect 1265 2370 1270 2410
rect 1335 2370 1340 2410
rect 1265 2365 1340 2370
rect 1385 2340 1415 3450
rect 1835 3060 1865 3450
rect 1835 2415 1865 3030
rect 1805 2410 1880 2415
rect 1805 2370 1810 2410
rect 1875 2370 1880 2410
rect 1805 2365 1880 2370
rect 1925 2340 1955 3450
rect 2375 3060 2405 3450
rect 2375 2415 2405 3030
rect 2345 2410 2420 2415
rect 2345 2370 2350 2410
rect 2415 2370 2420 2410
rect 2345 2365 2420 2370
rect 2465 2340 2495 3450
rect 2915 3060 2945 3450
rect 2915 2415 2945 3030
rect 2885 2410 2960 2415
rect 2885 2370 2890 2410
rect 2955 2370 2960 2410
rect 2885 2365 2960 2370
rect 3005 2340 3035 3450
rect 280 2335 355 2340
rect 280 2295 285 2335
rect 350 2295 355 2335
rect 280 2290 355 2295
rect 820 2335 895 2340
rect 820 2295 825 2335
rect 890 2295 895 2335
rect 820 2290 895 2295
rect 1360 2335 1435 2340
rect 1360 2295 1365 2335
rect 1430 2295 1435 2335
rect 1360 2290 1435 2295
rect 1900 2335 1975 2340
rect 1900 2295 1905 2335
rect 1970 2295 1975 2335
rect 1900 2290 1975 2295
rect 2440 2335 2515 2340
rect 2440 2295 2445 2335
rect 2510 2295 2515 2335
rect 2440 2290 2515 2295
rect 2980 2335 3055 2340
rect 2980 2295 2985 2335
rect 3050 2295 3055 2335
rect 2980 2290 3055 2295
rect 280 -7065 355 -7060
rect 280 -7105 285 -7065
rect 350 -7105 355 -7065
rect 280 -7110 355 -7105
rect 820 -7065 895 -7060
rect 820 -7105 825 -7065
rect 890 -7105 895 -7065
rect 820 -7110 895 -7105
rect 1360 -7065 1435 -7060
rect 1360 -7105 1365 -7065
rect 1430 -7105 1435 -7065
rect 1360 -7110 1435 -7105
rect 1900 -7065 1975 -7060
rect 1900 -7105 1905 -7065
rect 1970 -7105 1975 -7065
rect 1900 -7110 1975 -7105
rect 2440 -7065 2515 -7060
rect 2440 -7105 2445 -7065
rect 2510 -7105 2515 -7065
rect 2440 -7110 2515 -7105
rect 2980 -7065 3055 -7060
rect 2980 -7105 2985 -7065
rect 3050 -7105 3055 -7065
rect 2980 -7110 3055 -7105
rect 3425 -7065 3500 -7060
rect 3425 -7105 3430 -7065
rect 3495 -7095 4340 -7065
rect 3495 -7105 3500 -7095
rect 3425 -7110 3500 -7105
rect 185 -7140 260 -7135
rect 185 -7180 190 -7140
rect 255 -7180 260 -7140
rect 185 -7185 260 -7180
rect 215 -8220 245 -7185
rect 300 -8220 330 -7110
rect 725 -7140 800 -7135
rect 725 -7180 730 -7140
rect 795 -7180 800 -7140
rect 725 -7185 800 -7180
rect 755 -8220 785 -7185
rect 840 -8220 870 -7110
rect 1265 -7140 1340 -7135
rect 1265 -7180 1270 -7140
rect 1335 -7180 1340 -7140
rect 1265 -7185 1340 -7180
rect 1295 -8220 1325 -7185
rect 1380 -8220 1410 -7110
rect 1805 -7140 1880 -7135
rect 1805 -7180 1810 -7140
rect 1875 -7180 1880 -7140
rect 1805 -7185 1880 -7180
rect 1835 -8220 1865 -7185
rect 1920 -8220 1950 -7110
rect 2345 -7140 2420 -7135
rect 2345 -7180 2350 -7140
rect 2415 -7180 2420 -7140
rect 2345 -7185 2420 -7180
rect 2375 -8220 2405 -7185
rect 2460 -8220 2490 -7110
rect 2885 -7140 2960 -7135
rect 2885 -7180 2890 -7140
rect 2955 -7180 2960 -7140
rect 2885 -7185 2960 -7180
rect 2915 -8220 2945 -7185
rect 3000 -8220 3030 -7110
rect 170 -8225 255 -8220
rect 170 -8315 210 -8225
rect 250 -8315 255 -8225
rect 170 -8320 255 -8315
rect 290 -8225 375 -8220
rect 290 -8315 295 -8225
rect 335 -8315 375 -8225
rect 290 -8320 375 -8315
rect 170 -8595 205 -8320
rect 340 -8595 375 -8320
rect 710 -8225 795 -8220
rect 710 -8315 750 -8225
rect 790 -8315 795 -8225
rect 710 -8320 795 -8315
rect 830 -8225 915 -8220
rect 830 -8315 835 -8225
rect 875 -8315 915 -8225
rect 830 -8320 915 -8315
rect 710 -8595 745 -8320
rect 880 -8595 915 -8320
rect 1250 -8225 1335 -8220
rect 1250 -8315 1290 -8225
rect 1330 -8315 1335 -8225
rect 1250 -8320 1335 -8315
rect 1370 -8225 1455 -8220
rect 1370 -8315 1375 -8225
rect 1415 -8315 1455 -8225
rect 1370 -8320 1455 -8315
rect 1250 -8595 1285 -8320
rect 1420 -8595 1455 -8320
rect 1790 -8225 1875 -8220
rect 1790 -8315 1830 -8225
rect 1870 -8315 1875 -8225
rect 1790 -8320 1875 -8315
rect 1910 -8225 1995 -8220
rect 1910 -8315 1915 -8225
rect 1955 -8315 1995 -8225
rect 1910 -8320 1995 -8315
rect 1790 -8595 1825 -8320
rect 1960 -8595 1995 -8320
rect 2330 -8225 2415 -8220
rect 2330 -8315 2370 -8225
rect 2410 -8315 2415 -8225
rect 2330 -8320 2415 -8315
rect 2450 -8225 2535 -8220
rect 2450 -8315 2455 -8225
rect 2495 -8315 2535 -8225
rect 2450 -8320 2535 -8315
rect 2330 -8595 2365 -8320
rect 2500 -8595 2535 -8320
rect 2870 -8225 2955 -8220
rect 2870 -8315 2910 -8225
rect 2950 -8315 2955 -8225
rect 2870 -8320 2955 -8315
rect 2990 -8225 3075 -8220
rect 2990 -8315 2995 -8225
rect 3035 -8315 3075 -8225
rect 2990 -8320 3075 -8315
rect 2870 -8595 2905 -8320
rect 3040 -8595 3075 -8320
<< end >>
