* SPICE3 file created from pcbc.ext - technology: sky130A

X0 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X1 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X2 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X3 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X4 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X5 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X6 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X7 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X8 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X9 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X10 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X11 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X12 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X13 VP Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X14 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X15 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X16 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.6 as=0.5 ps=3.6 w=1 l=1
X17 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X18 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X19 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X20 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X21 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X22 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X23 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X24 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X25 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X26 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X27 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X28 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X29 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X30 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X31 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X32 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X33 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X34 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X35 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X36 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X37 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X38 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X39 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.6 as=0.2 ps=1.4 w=1 l=1
X40 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X41 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X42 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X43 Vdssat VP VP VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.56 ps=4.4 w=1 l=1
X44 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X45 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X46 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.6 as=0.5 ps=3.6 w=1 l=1
X47 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X48 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X49 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X50 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X51 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X52 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X53 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X54 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X55 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X56 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X57 Vdssat Vc Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X58 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X59 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X60 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X61 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X62 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X63 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X64 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X65 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X66 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X67 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X68 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X69 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X70 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X71 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X72 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X73 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X74 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X75 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X76 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X77 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.5 ps=3.6 w=1 l=1
X78 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X79 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X80 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X81 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X82 VP VP Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.56 pd=4.4 as=0.2 ps=1.4 w=1 l=1
X83 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X84 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X85 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X86 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X87 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X88 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X89 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X90 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X91 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X92 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X93 VP Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X94 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X95 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X96 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X97 Vdssat Vbg VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X98 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X99 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X100 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X101 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X102 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X103 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X104 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X105 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X106 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X107 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X108 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X109 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X110 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X111 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X112 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X113 Vdssat Vbg VP VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X114 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X115 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X116 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.6 as=0.2 ps=1.4 w=1 l=1
X117 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X118 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X119 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X120 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X121 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X122 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.5 ps=3.6 w=1 l=1
X123 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X124 VP VP Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.56 pd=4.4 as=0.2 ps=1.4 w=1 l=1
X125 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X126 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X127 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X128 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X129 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X130 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X131 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X132 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X133 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X134 Vdssat Vc Vc VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X135 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X136 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X137 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X138 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X139 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X140 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X141 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X142 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X143 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X144 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X145 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.6 as=0.5 ps=3.6 w=1 l=1
X146 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X147 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X148 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X149 Vc Vc Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X150 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X151 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X152 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X153 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X154 VN Vbn Vbg VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=0.4 ps=2.8 w=1 l=1
X155 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X156 Vbg Vbg Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X157 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X158 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.6 as=0.5 ps=3.6 w=1 l=1
X159 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X160 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X161 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X162 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X163 VN Vbn Vc VN sky130_fd_pr__nfet_01v8 ad=0.43 pd=3.1 as=3.58665 ps=25.33 w=1 l=10
X164 Vdssat Vbg Vbg VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=1
X165 Vc Vbn VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.43 ps=3.1 w=1 l=10
X166 Vc VN VN VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=10
X167 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X168 VN VN Vc VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=10
X169 Vc Vc Vdssat VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X170 Vbg Vbn VN VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.43 ps=3.1 w=1 l=1
X171 Vdssat VP VP VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.56 ps=4.4 w=1 l=1
.end

