magic
tech sky130A
timestamp 1762200811
<< nwell >>
rect -90 250 200 490
<< nmos >>
rect 0 0 50 200
rect 90 0 140 200
<< pmos >>
rect 0 270 50 470
rect 90 270 140 470
<< ndiff >>
rect -40 110 0 200
rect -40 90 -30 110
rect -10 90 0 110
rect -40 0 0 90
rect 50 190 90 200
rect 50 170 60 190
rect 80 170 90 190
rect 50 0 90 170
rect 140 110 180 200
rect 140 90 150 110
rect 170 90 180 110
rect 140 0 180 90
<< pdiff >>
rect -40 380 0 470
rect -40 360 -30 380
rect -10 360 0 380
rect -40 270 0 360
rect 50 460 90 470
rect 50 440 60 460
rect 80 440 90 460
rect 50 300 90 440
rect 50 280 60 300
rect 80 280 90 300
rect 50 270 90 280
rect 140 380 180 470
rect 140 360 150 380
rect 170 360 180 380
rect 140 270 180 360
<< ndiffc >>
rect -30 90 -10 110
rect 60 170 80 190
rect 150 90 170 110
<< pdiffc >>
rect -30 360 -10 380
rect 60 440 80 460
rect 60 280 80 300
rect 150 360 170 380
<< psubdiff >>
rect -70 110 -40 200
rect -50 90 -40 110
rect -70 0 -40 90
<< nsubdiff >>
rect -70 380 -40 470
rect -50 360 -40 380
rect -70 270 -40 360
<< psubdiffcont >>
rect -70 90 -50 110
<< nsubdiffcont >>
rect -70 360 -50 380
<< poly >>
rect 0 470 50 490
rect 90 470 140 490
rect 0 250 50 270
rect 90 250 140 270
rect 10 220 40 250
rect 100 220 130 250
rect 0 200 50 220
rect 90 200 140 220
rect 0 -10 50 0
rect 90 -10 140 0
rect 0 -20 140 -10
rect 0 -40 60 -20
rect 80 -40 140 -20
rect 0 -50 140 -40
<< polycont >>
rect 60 -40 80 -20
<< locali >>
rect 50 460 90 490
rect 50 440 60 460
rect 80 440 90 460
rect 50 430 90 440
rect -70 380 180 390
rect -50 360 -30 380
rect -10 360 150 380
rect 170 360 180 380
rect -70 350 180 360
rect 50 300 90 310
rect 50 280 60 300
rect 80 280 90 300
rect 50 190 90 280
rect 50 170 60 190
rect 80 170 90 190
rect 50 160 90 170
rect -70 110 180 120
rect -50 90 -30 110
rect -10 90 150 110
rect 170 90 180 110
rect -70 80 180 90
rect -70 -20 90 -10
rect -70 -40 60 -20
rect 80 -40 90 -20
rect -70 -50 90 -40
<< labels >>
rlabel locali -70 -30 -70 -30 7 A
port 1 w
rlabel locali 70 490 70 490 1 Y
port 2 n
rlabel nsubdiffcont -70 370 -70 370 7 VP
port 3 w
rlabel psubdiffcont -70 100 -70 100 7 VN
port 4 w
<< end >>
