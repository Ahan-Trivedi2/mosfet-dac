* SPICE3 file created from full.ext - technology: sky130A

X0 dac_0/a_6220_2110# inv_0/A dac_0/a_6220_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X1 dac_0/a_2270_n1450# inv_7/VP dac_0/a_2270_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X2 dac_0/a_3350_n7120# inv_7/VP dac_0/a_3350_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X3 dac_0/a_1900_3210# inv_7/A dac_0/a_1900_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X4 dac_0/a_4060_n7120# inv_7/VP dac_0/a_4060_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X5 inv_7/VN inv_7/VN fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X6 dac_0/a_110_n350# inv_7/VP dac_0/a_110_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X7 inv_7/VN inv_7/VN dac_0/a_3350_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X8 dac_0/a_3350_n2550# inv_7/VP dac_0/a_2270_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X9 inv_7/VN inv_7/VN dac_0/a_4430_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X10 dac_0/a_4060_n2550# inv_7/VP dac_0/a_3350_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X11 dac_0/a_4430_n8220# inv_7/VP dac_0/a_4430_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X12 dac_0/a_5140_n8220# inv_7/VP dac_0/a_5140_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X13 dac_0/a_5140_4310# inv_1/A dac_0/a_5140_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X14 dac_0/a_4060_n10730# inv_2/A dac_0/a_4060_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X15 dac_0/a_4430_3210# inv_2/Y dac_0/a_4430_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X16 dac_0/a_3350_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X17 dac_0/a_n260_n9320# inv_7/VP dac_0/a_n260_n10730# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X18 dac_0/a_4430_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X19 inv_7/VN inv_7/VN dac_0/a_110_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X20 dac_0/a_1190_n10420# inv_7/VP dac_0/a_1900_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X21 dac_0/a_4060_n14030# inv_2/A fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X22 dac_0/a_5140_n11830# inv_1/A dac_0/a_5140_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X23 dac_0/a_6220_n10730# inv_0/Y dac_0/a_6590_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X24 inv_7/VN inv_7/VN fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X25 inv_7/VN inv_7/VN fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X26 dac_0/a_820_n8220# inv_7/VP dac_0/a_820_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X27 fvf_1/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X28 dac_0/a_2270_n9320# inv_7/VP dac_0/a_2270_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X29 dac_0/a_4430_n350# inv_7/VP dac_0/a_4430_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X30 dac_0/a_1900_n1450# inv_7/VP dac_0/a_1900_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X31 dac_0/a_6590_n14030# inv_0/Y fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X32 dac_0/a_6220_n12930# inv_0/A dac_0/a_6220_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X33 inv_7/VN inv_7/VN fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X34 dac_0/a_5140_n350# inv_7/VP dac_0/a_5140_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X35 dac_0/a_2270_n10420# inv_7/VP dac_0/a_2980_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X36 dac_0/a_4430_n10420# inv_7/VP dac_0/a_5510_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X37 dac_0/a_1900_n12930# inv_7/A dac_0/a_1900_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X38 fvf_0/Vin inv_3/Y dac_0/a_3350_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X39 dac_0/a_3350_750# inv_7/VP dac_0/a_3350_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X40 dac_0/a_110_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X41 dac_0/a_5510_n10420# inv_7/VP dac_0/a_6220_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X42 dac_0/a_110_3210# inv_4/Y dac_0/a_110_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X43 dac_0/a_820_3210# inv_6/A dac_0/a_820_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X44 dac_0/a_2980_n1450# inv_7/VP dac_0/a_2980_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X45 dac_0/a_5510_n1450# inv_7/VP dac_0/a_5510_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X46 dac_0/a_4060_3210# inv_2/A dac_0/a_4060_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X47 dac_0/a_6220_n1450# inv_7/VP dac_0/a_6220_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X48 dac_0/a_5510_n10420# inv_7/VP dac_0/a_6590_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X49 dac_0/a_7300_n7120# inv_7/VP dac_0/a_7300_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X50 dac_0/a_3350_2110# inv_3/Y dac_0/a_2980_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X51 dac_0/a_820_n350# inv_7/VP dac_0/a_820_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X52 dac_0/a_n260_n11830# inv_4/A dac_0/a_n260_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X53 fvf_0/Vin inv_0/Y dac_0/a_6590_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X54 dac_0/a_6590_750# inv_7/VP dac_0/a_6590_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X55 dac_0/a_820_n10730# inv_6/Y dac_0/a_1190_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X56 dac_0/a_6590_n1450# inv_7/VP dac_0/a_6590_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X57 dac_0/a_7300_n2550# inv_7/VP dac_0/a_6590_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X58 fvf_1/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X59 dac_0/a_1190_n14030# inv_6/Y fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X60 dac_0/a_2270_n11830# inv_7/Y dac_0/a_2270_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X61 dac_0/a_6590_2110# inv_0/Y dac_0/a_6220_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X62 inv_7/VN inv_7/VN dac_0/Iin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X63 dac_0/a_5510_n9320# inv_7/VP dac_0/a_5510_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X64 dac_0/a_2270_4310# inv_7/Y dac_0/a_2270_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X65 dac_0/a_2980_4310# inv_3/A dac_0/a_2980_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X66 fvf_0/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X67 dac_0/a_3350_n12930# inv_3/Y dac_0/a_3350_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X68 dac_0/a_n260_n8220# inv_7/VP dac_0/a_n260_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X69 dac_0/a_110_n12930# inv_4/Y dac_0/a_110_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X70 dac_0/Iin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X71 inv_7/VN inv_7/VN fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X72 dac_0/a_4060_n10730# inv_2/Y dac_0/a_4430_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X73 dac_0/a_820_n9320# inv_7/VP dac_0/a_820_n10730# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X74 fvf_0/Vin inv_7/VP dac_0/a_7300_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X75 inv_7/VN inv_7/VN fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X76 dac_0/a_n260_n350# inv_7/VP dac_0/a_n260_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X77 dac_0/a_4430_n14030# inv_2/Y fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X78 dac_0/a_5510_n11830# inv_1/Y dac_0/a_5510_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X79 dac_0/a_1190_3210# inv_6/Y dac_0/a_1190_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X80 dac_0/a_1190_n7120# inv_7/VP dac_0/a_1190_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X81 dac_0/a_2980_n10730# inv_3/A dac_0/a_2980_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X82 inv_7/VN inv_7/VN dac_0/a_1190_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X83 fvf_0/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X84 dac_0/a_n260_3210# inv_4/A dac_0/a_n260_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X85 dac_0/a_2980_n14030# inv_3/A fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X86 inv_7/VN inv_7/VN fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X87 dac_0/a_1190_n2550# inv_7/VP dac_0/a_110_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X88 dac_0/a_2270_n8220# inv_7/VP dac_0/a_2270_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X89 dac_0/a_110_n7120# inv_7/VP dac_0/a_110_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X90 dac_0/a_820_n11830# inv_6/A dac_0/a_820_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X91 dac_0/a_6220_4310# inv_0/A dac_0/a_6220_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X92 dac_0/a_5510_3210# inv_1/Y dac_0/a_5510_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X93 dac_0/a_1190_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X94 fvf_1/Vin inv_7/A dac_0/a_1900_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X95 dac_0/a_1900_750# inv_7/VP dac_0/a_1900_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X96 dac_0/a_110_n2550# inv_7/VP dac_0/Iin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X97 fvf_1/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X98 dac_0/a_2270_n350# inv_7/VP dac_0/a_2270_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X99 dac_0/a_2270_n10420# inv_7/VP dac_0/a_3350_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X100 dac_0/a_1900_2110# inv_7/A dac_0/a_1900_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X101 dac_0/a_3350_n10420# inv_7/VP dac_0/a_4060_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X102 dac_0/a_6220_n9320# inv_7/VP dac_0/a_6220_n10730# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X103 inv_7/VN inv_7/VN fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X104 fvf_0/Vin inv_2/Y dac_0/a_4430_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X105 inv_7/VN inv_7/VN dac_0/a_1190_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X106 dac_0/a_4060_n12930# inv_2/A dac_0/a_4060_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X107 dac_0/a_1900_n9320# inv_7/VP dac_0/a_1900_n10730# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X108 dac_0/a_4430_750# inv_7/VP dac_0/a_4430_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X109 dac_0/a_3350_n1450# inv_7/VP dac_0/a_3350_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X110 dac_0/a_4060_n1450# inv_7/VP dac_0/a_4060_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X111 dac_0/a_4430_n7120# inv_7/VP dac_0/a_4430_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X112 dac_0/a_1900_n8220# inv_7/VP dac_0/a_1900_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X113 dac_0/a_5140_n7120# inv_7/VP dac_0/a_5140_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X114 dac_0/a_6590_n12930# inv_0/Y dac_0/a_6590_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X115 dac_0/a_5140_3210# inv_1/A dac_0/a_5140_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X116 inv_7/VN inv_7/VN dac_0/a_2270_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X117 inv_7/VN inv_7/VN dac_0/a_4430_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X118 inv_7/VN inv_7/VN dac_0/a_5510_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X119 dac_0/a_4430_2110# inv_2/Y dac_0/a_4060_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X120 dac_0/a_4430_n2550# inv_7/VP dac_0/a_3350_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X121 dac_0/a_1190_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X122 dac_0/a_5140_n2550# inv_7/VP dac_0/a_4430_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X123 dac_0/a_5140_n10730# inv_1/A dac_0/a_5140_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X124 dac_0/a_5510_n8220# inv_7/VP dac_0/a_5510_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X125 dac_0/a_2980_n8220# inv_7/VP dac_0/a_2980_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X126 dac_0/a_6220_n8220# inv_7/VP dac_0/a_6220_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X127 fvf_0/Vin inv_4/Y dac_0/a_110_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X128 fvf_1/Vin inv_6/A dac_0/a_820_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X129 dac_0/a_110_750# inv_7/VP dac_0/a_110_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X130 dac_0/a_820_750# inv_7/VP dac_0/a_820_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X131 inv_7/VN inv_7/VN dac_0/a_5510_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X132 dac_0/a_820_n7120# inv_7/VP dac_0/a_820_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X133 dac_0/a_1900_n350# inv_7/VP dac_0/a_1900_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X134 dac_0/a_2270_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X135 dac_0/a_4430_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X136 dac_0/a_5140_n14030# inv_1/A fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X137 dac_0/a_6220_n11830# inv_0/A dac_0/a_6220_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X138 fvf_1/Vin inv_2/A dac_0/a_4060_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X139 dac_0/a_4060_750# inv_7/VP dac_0/a_4060_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X140 dac_0/a_5510_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X141 dac_0/a_1900_n11830# inv_7/A dac_0/a_1900_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X142 dac_0/a_6590_n8220# inv_7/VP dac_0/a_6590_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X143 dac_0/a_3350_4310# inv_3/Y dac_0/a_3350_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X144 dac_0/a_820_n2550# inv_7/VP dac_0/a_110_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X145 fvf_1/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X146 dac_0/a_3350_n9320# inv_7/VP dac_0/a_3350_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X147 dac_0/a_110_2110# inv_4/Y dac_0/a_n260_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X148 dac_0/a_820_2110# inv_6/A dac_0/a_820_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X149 fvf_1/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X150 dac_0/a_1190_n12930# inv_6/Y dac_0/a_1190_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X151 dac_0/a_2980_n350# inv_7/VP dac_0/a_2980_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X152 dac_0/a_5510_n350# inv_7/VP dac_0/a_5510_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X153 dac_0/a_5510_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X154 dac_0/a_4060_2110# inv_2/A dac_0/a_4060_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X155 dac_0/a_6220_n350# inv_7/VP dac_0/a_6220_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X156 dac_0/a_110_n9320# inv_7/VP dac_0/a_110_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X157 dac_0/a_6590_n10420# inv_7/VP dac_0/a_7300_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X158 dac_0/a_n260_n10730# inv_4/A dac_0/a_n260_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X159 dac_0/a_6590_4310# inv_0/Y dac_0/a_6590_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X160 inv_7/VN inv_7/VN fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X161 inv_7/VN inv_7/VN fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X162 dac_0/a_6590_n350# inv_7/VP dac_0/a_6590_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X163 dac_0/a_7300_n1450# inv_7/VP dac_0/a_7300_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X164 dac_0/a_n260_n14030# inv_4/A fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X165 dac_0/a_1900_n10730# inv_7/Y dac_0/a_2270_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X166 dac_0/a_2270_3210# inv_7/Y dac_0/a_2270_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X167 dac_0/a_2980_3210# inv_3/A dac_0/a_2980_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X168 dac_0/a_2270_n14030# inv_7/Y fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X169 dac_0/a_3350_n11830# inv_3/Y dac_0/a_3350_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X170 dac_0/a_n260_n7120# inv_7/VP dac_0/a_n260_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X171 fvf_0/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X172 dac_0/a_4430_n12930# inv_2/Y dac_0/a_4430_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X173 dac_0/a_110_n11830# inv_4/Y dac_0/a_110_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X174 dac_0/a_n260_n2550# inv_7/VP dac_0/Iin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X175 fvf_0/Vin inv_6/Y dac_0/a_1190_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X176 dac_0/a_1190_750# inv_7/VP dac_0/a_1190_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X177 fvf_0/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X178 dac_0/a_2980_n12930# inv_3/A dac_0/a_2980_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X179 fvf_1/Vin inv_4/A dac_0/a_n260_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X180 dac_0/a_n260_750# inv_7/VP dac_0/a_n260_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X181 dac_0/a_5140_n10730# inv_1/Y dac_0/a_5510_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X182 dac_0/a_1190_2110# inv_6/Y dac_0/a_820_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X183 dac_0/a_110_n10420# inv_7/VP dac_0/a_1190_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X184 dac_0/a_5510_n14030# inv_1/Y fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X185 dac_0/a_n260_2110# inv_4/A dac_0/a_n260_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X186 inv_7/VN inv_7/VN fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X187 fvf_0/Vin inv_1/Y dac_0/a_5510_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X188 dac_0/a_1190_n1450# inv_7/VP dac_0/a_1190_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X189 dac_0/a_4060_n9320# inv_7/VP dac_0/a_4060_n10730# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X190 dac_0/a_5510_750# inv_7/VP dac_0/a_5510_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X191 dac_0/a_2270_n7120# inv_7/VP dac_0/a_2270_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X192 inv_7/VN inv_7/VN dac_0/a_2270_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X193 dac_0/a_6590_n9320# inv_7/VP dac_0/a_6590_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X194 inv_7/VN inv_7/VN dac_0/a_3350_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X195 dac_0/Iin inv_7/VP dac_0/a_110_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X196 dac_0/a_820_n10730# inv_6/A dac_0/a_820_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X197 dac_0/a_6220_3210# inv_0/A dac_0/a_6220_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X198 dac_0/a_5510_2110# inv_1/Y dac_0/a_5140_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X199 dac_0/a_2270_n2550# inv_7/VP dac_0/a_1190_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X200 dac_0/a_3350_n8220# inv_7/VP dac_0/a_3350_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X201 dac_0/a_1900_4310# inv_7/A dac_0/a_1900_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X202 dac_0/a_820_n14030# inv_6/A fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X203 dac_0/a_4060_n8220# inv_7/VP dac_0/a_4060_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X204 dac_0/a_110_n1450# inv_7/VP dac_0/a_110_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X205 dac_0/a_2270_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X206 dac_0/a_3350_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X207 fvf_1/Vin inv_1/A dac_0/a_5140_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X208 dac_0/a_5140_750# inv_7/VP dac_0/a_5140_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X209 dac_0/a_4060_n11830# inv_2/A dac_0/a_4060_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X210 dac_0/a_4430_4310# inv_2/Y dac_0/a_4430_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X211 dac_0/a_7300_n9320# inv_7/VP fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X212 dac_0/a_3350_n350# inv_7/VP dac_0/a_3350_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X213 dac_0/a_4060_n350# inv_7/VP dac_0/a_4060_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X214 dac_0/a_3350_n10420# inv_7/VP dac_0/a_4430_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X215 dac_0/a_1900_n7120# inv_7/VP dac_0/a_1900_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X216 fvf_1/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X217 dac_0/a_5140_n12930# inv_1/A dac_0/a_5140_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X218 dac_0/a_1190_n9320# inv_7/VP dac_0/a_1190_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X219 dac_0/a_4430_n10420# inv_7/VP dac_0/a_5140_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X220 dac_0/a_6590_n11830# inv_0/Y dac_0/a_6590_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X221 dac_0/a_5140_2110# inv_1/A dac_0/a_5140_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X222 dac_0/a_4430_n1450# inv_7/VP dac_0/a_4430_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X223 dac_0/a_1900_n2550# inv_7/VP dac_0/a_1190_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X224 fvf_0/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X225 dac_0/a_5140_n1450# inv_7/VP dac_0/a_5140_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X226 dac_0/a_2980_n7120# inv_7/VP dac_0/a_2980_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X227 dac_0/a_5510_n7120# inv_7/VP dac_0/a_5510_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X228 inv_7/VN inv_7/VN fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X229 dac_0/a_6220_n7120# inv_7/VP dac_0/a_6220_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X230 dac_0/a_110_4310# inv_4/Y dac_0/a_110_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X231 dac_0/a_820_4310# inv_6/A dac_0/a_820_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X232 inv_7/VN inv_7/VN dac_0/a_6590_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X233 dac_0/a_110_n10420# inv_7/VP dac_0/a_820_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X234 dac_0/a_2980_n2550# inv_7/VP dac_0/a_2270_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X235 dac_0/a_5510_n2550# inv_7/VP dac_0/a_4430_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X236 dac_0/a_6220_n10730# inv_0/A dac_0/a_6220_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X237 dac_0/a_4060_4310# inv_2/A dac_0/a_4060_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X238 dac_0/a_6220_n2550# inv_7/VP dac_0/a_5510_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X239 dac_0/a_6590_n7120# inv_7/VP dac_0/a_6590_n8220# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X240 dac_0/a_1900_n10730# inv_7/A dac_0/a_1900_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X241 dac_0/a_7300_n8220# inv_7/VP dac_0/a_7300_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X242 dac_0/a_3350_3210# inv_3/Y dac_0/a_3350_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X243 dac_0/a_820_n1450# inv_7/VP dac_0/a_820_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X244 dac_0/a_6220_n14030# inv_0/A fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X245 dac_0/a_n260_n12930# inv_4/A dac_0/a_n260_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X246 inv_7/VN inv_7/VN fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X247 dac_0/a_1900_n14030# inv_7/A fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X248 dac_0/a_1190_n11830# inv_6/Y dac_0/a_1190_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X249 dac_0/a_6590_n2550# inv_7/VP dac_0/a_5510_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X250 dac_0/a_6590_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X251 dac_0/a_4430_n9320# inv_7/VP dac_0/a_4430_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X252 fvf_0/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X253 dac_0/a_2270_n12930# inv_7/Y dac_0/a_2270_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X254 dac_0/a_6590_3210# inv_0/Y dac_0/a_6590_2110# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X255 dac_0/a_2980_n9320# inv_7/VP dac_0/a_2980_n10730# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X256 fvf_0/Vin inv_7/Y dac_0/a_2270_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X257 fvf_1/Vin inv_3/A dac_0/a_2980_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X258 dac_0/a_2270_750# inv_7/VP dac_0/a_2270_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X259 dac_0/a_2980_750# inv_7/VP dac_0/a_2980_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X260 dac_0/a_7300_n350# inv_7/VP dac_0/a_7300_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X261 dac_0/a_2270_2110# inv_7/Y dac_0/a_1900_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X262 dac_0/a_2980_2110# inv_3/A dac_0/a_2980_750# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X263 dac_0/a_2980_n10730# inv_3/Y dac_0/a_3350_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X264 dac_0/Iin inv_7/VP dac_0/a_n260_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X265 dac_0/a_3350_n14030# inv_3/Y fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X266 dac_0/a_4430_n11830# inv_2/Y dac_0/a_4430_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X267 inv_7/VN inv_7/VN dac_0/a_110_n10420# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X268 fvf_0/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X269 dac_0/a_n260_n10730# inv_4/Y dac_0/a_110_n11830# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X270 dac_0/a_n260_n1450# inv_7/VP dac_0/a_n260_n2550# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X271 dac_0/a_5510_n12930# inv_1/Y dac_0/a_5510_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X272 dac_0/a_1190_4310# inv_6/Y dac_0/a_1190_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X273 dac_0/a_1190_n8220# inv_7/VP dac_0/a_1190_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X274 dac_0/a_110_n14030# inv_4/Y fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X275 dac_0/a_2980_n11830# inv_3/A dac_0/a_2980_n12930# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X276 dac_0/a_n260_4310# inv_4/A dac_0/a_n260_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X277 fvf_1/Vin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X278 dac_0/a_110_750# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X279 inv_7/VN inv_7/VN dac_0/Iin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X280 dac_0/a_110_n8220# inv_7/VP dac_0/a_110_n9320# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X281 dac_0/a_820_n12930# inv_6/A dac_0/a_820_n14030# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X282 fvf_1/Vin inv_0/A dac_0/a_6220_4310# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X283 dac_0/a_5510_4310# inv_1/Y dac_0/a_5510_3210# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X284 dac_0/a_6220_750# inv_7/VP dac_0/a_6220_n350# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X285 dac_0/a_1190_n350# inv_7/VP dac_0/a_1190_n1450# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X286 inv_7/VN inv_7/VN fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.375 pd=2.5 as=0.1875 ps=1.25 w=0.75 l=5
X287 dac_0/Iin inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X288 dac_0/a_1190_n10420# inv_7/VP dac_0/a_2270_n7120# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.1875 ps=1.25 w=0.75 l=5
X289 dac_0/a_5140_n9320# inv_7/VP dac_0/a_5140_n10730# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.1875 pd=1.25 as=0.375 ps=2.5 w=0.75 l=5
X290 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X291 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X292 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X293 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X294 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X295 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X296 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X297 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X298 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X299 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X300 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X301 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X302 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X303 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X304 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X305 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X306 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X307 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X308 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X309 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X310 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X311 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X312 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X313 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X314 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X315 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X316 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X317 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X318 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X319 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X320 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X321 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X322 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X323 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X324 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X325 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X326 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X327 fvf_1/VP pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X328 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X329 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X330 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X331 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X332 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X333 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X334 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X335 pcbc_0/Vc pcbc_0/Vc pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X336 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X337 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X338 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X339 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X340 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X341 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X342 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X343 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X344 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X345 pcbc_0/Vc pcbc_0/Vc pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X346 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X347 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X348 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X349 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X350 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X351 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X352 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X353 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X354 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X355 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X356 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X357 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X358 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X359 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X360 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X361 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X362 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X363 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X364 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X365 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X366 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X367 pcbc_0/a_8360_6840# pcbc_0/Vc pcbc_0/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X368 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X369 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X370 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X371 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X372 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X373 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X374 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X375 fvf_1/VP fvf_1/VP pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X376 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X377 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X378 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X379 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X380 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X381 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X382 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X383 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X384 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X385 fvf_1/VP fvf_1/VP pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X386 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X387 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X388 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X389 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X390 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X391 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X392 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X393 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X394 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X395 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X396 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X397 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X398 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X399 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X400 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X401 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X402 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X403 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X404 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X405 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X406 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X407 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X408 pcbc_0/a_8360_6840# fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X409 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X410 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X411 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X412 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X413 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X414 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X415 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X416 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X417 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X418 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X419 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X420 fvf_1/VP pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X421 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X422 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X423 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X424 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X425 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X426 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X427 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X428 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X429 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X430 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X431 pcbc_0/a_8360_6840# fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X432 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X433 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X434 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X435 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X436 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X437 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X438 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X439 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X440 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X441 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X442 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X443 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X444 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X445 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X446 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X447 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X448 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X449 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X450 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X451 inv_7/VN bbg_0/VBN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X452 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X453 pcbc_0/Vc inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X454 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X455 inv_7/VN inv_7/VN pcbc_0/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X456 pcbc_0/a_8360_6840# pcbc_0/Vc pcbc_0/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X457 pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# pcbc_0/a_8360_6840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X458 pcbc_0/a_8360_6840# pcbc_0/a_8320_6920# pcbc_0/a_8320_6920# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X459 pcbc_0/Vc bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X460 inv_7/VN bbg_0/VBN pcbc_0/a_8320_6920# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X461 pcbc_0/a_8320_6920# bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X462 fvf_1/VP ccm_0/a_3280_100# ccm_0/a_3480_1180# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X463 ccm_0/a_3280_100# fvf_1/Vc ccm_0/a_2200_100# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.87 pd=5.3 as=0.58 ps=3.53 w=2 l=5
X464 ccm_0/a_2200_100# Vcn inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.58 pd=3.53 as=2.14 ps=7 w=2 l=5
X465 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=108.96002 ps=551.005 w=2 l=5
X466 ccm_0/Vout fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=1.47 ps=5.9 w=2 l=5
X467 fvf_1/VP ccm_0/a_3280_100# ccm_0/a_3280_100# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.87 ps=5.3 w=2 l=5
X468 ccm_0/Vout fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=1.47 ps=5.9 w=2 l=5
X469 inv_7/VN Vcn ccm_0/a_n80_100# inv_7/VN sky130_fd_pr__nfet_01v8 ad=2.14 pd=7 as=0.58 ps=3.53 w=2 l=5
X470 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0 ps=0 w=2 l=5
X471 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0 ps=0 w=2 l=5
X472 ccm_0/Vout pcbc_0/Vc ccm_0/a_n1360_1180# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X473 ccm_0/Vout pcbc_0/Vc ccm_0/a_n1360_1180# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X474 fvf_1/VP fvf_1/VP ccm_0/Vout fvf_1/VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0.58 ps=3.53 w=2 l=5
X475 fvf_1/VP fvf_1/VP ccm_0/Vout fvf_1/VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0.58 ps=3.53 w=2 l=5
X476 ccm_0/a_2200_100# Vcn inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.58 pd=3.53 as=2.14 ps=7 w=2 l=5
X477 ccm_0/a_n80_100# fvf_1/Vc ccm_0/a_n2360_60# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.58 pd=3.53 as=0.87 ps=5.3 w=2 l=5
X478 inv_7/VN Vcn ccm_0/a_n80_100# inv_7/VN sky130_fd_pr__nfet_01v8 ad=2.14 pd=7 as=0.58 ps=3.53 w=2 l=5
X479 ccm_0/a_n1360_1180# ccm_0/a_n2360_60# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X480 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0 ps=0 w=2 l=5
X481 ccm_0/a_n1360_1180# ccm_0/a_n2360_60# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X482 ccm_0/a_n2360_60# ccm_0/a_n2360_60# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.87 pd=5.3 as=0.58 ps=3.53 w=2 l=5
X483 ccm_0/a_n80_100# fvf_1/Vc ccm_0/a_n2360_60# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.58 pd=3.53 as=0.87 ps=5.3 w=2 l=5
X484 ccm_0/a_3480_1180# pcbc_0/Vc ccm_0/Vout fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X485 ccm_0/a_3480_1180# pcbc_0/Vc ccm_0/Vout fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X486 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0 ps=0 w=2 l=5
X487 ccm_0/a_3280_100# fvf_1/Vc ccm_0/a_2200_100# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.87 pd=5.3 as=0.58 ps=3.53 w=2 l=5
X488 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0 ps=0 w=2 l=5
X489 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=1.47 pd=5.9 as=0 ps=0 w=2 l=5
X490 ccm_0/a_n2360_60# ccm_0/a_n2360_60# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.87 pd=5.3 as=0.58 ps=3.53 w=2 l=5
X491 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0 ps=0 w=2 l=5
X492 fvf_1/VP ccm_0/a_3280_100# ccm_0/a_3480_1180# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.58 ps=3.53 w=2 l=5
X493 fvf_1/VP ccm_0/a_3280_100# ccm_0/a_3280_100# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.58 pd=3.53 as=0.87 ps=5.3 w=2 l=5
X494 inv_0/Y inv_0/A inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.5
X495 inv_0/Y inv_0/A inv_7/VP inv_7/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.5
X496 inv_7/VP inv_0/A inv_0/Y inv_7/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5
X497 inv_7/VN inv_0/A inv_0/Y inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.5
X498 inv_1/Y inv_1/A inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=116.75 ps=631.40002 w=2 l=0.5
X499 inv_1/Y inv_1/A inv_7/VP inv_7/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=12.08 ps=74.8 w=2 l=0.5
X500 inv_7/VP inv_1/A inv_1/Y inv_7/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X501 inv_7/VN inv_1/A inv_1/Y inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X502 inv_2/Y inv_2/A inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X503 inv_2/Y inv_2/A inv_7/VP inv_7/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X504 inv_7/VP inv_2/A inv_2/Y inv_7/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X505 inv_7/VN inv_2/A inv_2/Y inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X506 inv_3/Y inv_3/A inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X507 inv_3/Y inv_3/A inv_7/VP inv_7/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X508 inv_7/VP inv_3/A inv_3/Y inv_7/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X509 inv_7/VN inv_3/A inv_3/Y inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X510 inv_4/Y inv_4/A inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X511 inv_4/Y inv_4/A inv_7/VP inv_7/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X512 inv_7/VP inv_4/A inv_4/Y inv_7/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X513 inv_7/VN inv_4/A inv_4/Y inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X514 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X515 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X516 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X517 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X518 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X519 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X520 ncbc_0/a_n560_3080# fvf_1/Vc fvf_1/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X521 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X522 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X523 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X524 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X525 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X526 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X527 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X528 fvf_1/Vc fvf_1/Vc ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X529 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X530 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X531 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X532 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X533 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X534 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X535 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X536 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X537 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X538 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X539 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X540 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X541 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X542 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X543 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X544 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X545 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X546 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X547 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X548 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X549 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X550 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X551 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X552 fvf_1/Vc fvf_1/Vc ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X553 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X554 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X555 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X556 ncbc_0/a_n560_3080# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X557 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X558 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X559 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X560 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X561 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X562 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X563 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X564 inv_7/VN ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X565 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X566 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X567 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X568 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X569 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X570 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X571 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X572 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X573 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X574 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X575 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X576 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X577 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X578 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X579 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X580 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X581 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X582 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X583 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X584 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X585 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X586 inv_7/VN inv_7/VN ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X587 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X588 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X589 ncbc_0/a_n560_3080# fvf_1/Vc fvf_1/Vc inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X590 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X591 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X592 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X593 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X594 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X595 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X596 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X597 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X598 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X599 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X600 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X601 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X602 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X603 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X604 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X605 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X606 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X607 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X608 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X609 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X610 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X611 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X612 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X613 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X614 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X615 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X616 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X617 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X618 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X619 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X620 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X621 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X622 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X623 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X624 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=2.69333 ps=14 w=10 l=1
X625 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X626 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X627 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X628 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X629 inv_7/VN ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=5
X630 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X631 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=5
X632 ncbc_0/a_n560_3080# inv_7/VN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=7.9 ps=22.1 w=10 l=1
X633 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X634 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X635 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X636 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X637 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X638 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X639 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X640 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X641 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=2.69333 pd=14 as=4.04 ps=21 w=10 l=1
X642 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X643 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X644 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X645 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X646 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X647 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X648 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X649 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X650 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X651 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X652 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X653 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X654 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X655 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X656 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X657 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X658 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X659 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X660 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X661 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X662 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X663 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X664 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X665 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X666 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X667 inv_7/VN inv_7/VN ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=7.9 pd=22.1 as=2.69333 ps=14 w=10 l=1
X668 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X669 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X670 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X671 ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# ncbc_0/a_n560_3080# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X672 fvf_1/VP fvf_1/VP fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=3.58665 ps=25.33 w=1 l=1
X673 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X674 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X675 fvf_1/VP fvf_1/Vbp ncbc_0/a_n600_3160# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X676 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X677 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X678 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X679 ncbc_0/a_n600_3160# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X680 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X681 fvf_1/VP fvf_1/Vbp fvf_1/Vc fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=3.58665 ps=25.33 w=1 l=1
X682 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X683 ncbc_0/a_n560_3080# ncbc_0/a_n600_3160# ncbc_0/a_n600_3160# inv_7/VN sky130_fd_pr__nfet_01v8 ad=4.04 pd=21 as=4.04 ps=21 w=10 l=1
X684 fvf_1/Vc fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.4 ps=2.8 w=1 l=1
X685 fvf_1/Vc fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=3.58665 pd=25.33 as=0.2 ps=1.4 w=1 l=1
X686 inv_7/Y inv_7/A inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X687 inv_7/Y inv_7/A inv_7/VP inv_7/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X688 inv_7/VP inv_7/A inv_7/Y inv_7/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X689 inv_7/VN inv_7/A inv_7/Y inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X690 inv_6/Y inv_6/A inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X691 inv_6/Y inv_6/A inv_7/VP inv_7/VP sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.5
X692 inv_7/VP inv_6/A inv_6/Y inv_7/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X693 inv_7/VN inv_6/A inv_6/Y inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X694 inv_7/VN bbg_0/a_460_n780# bbg_0/a_n200_n840# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X695 bbg_0/a_460_n780# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X696 bbg_0/a_460_n780# bbg_0/a_460_n780# bbg_0/RES inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X697 fvf_1/VP fvf_1/Vbp bbg_0/a_460_n780# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X698 bbg_0/a_n200_n840# bbg_0/a_460_n780# inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X699 fvf_1/VP bbg_0/a_n200_n840# bbg_0/a_n200_n840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X700 inv_7/VN bbg_0/VBN fvf_1/Vbp inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X701 fvf_1/Vbp bbg_0/a_n200_n840# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X702 bbg_0/VBN fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X703 bbg_0/a_n200_n840# bbg_0/a_460_n780# inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X704 bbg_0/RES bbg_0/a_460_n780# bbg_0/a_460_n780# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X705 fvf_1/VP fvf_1/Vbp bbg_0/VBN fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X706 fvf_1/VP fvf_1/Vbp bbg_0/VBN fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X707 fvf_1/Vbp bbg_0/a_n200_n840# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X708 bbg_0/a_n200_n840# bbg_0/a_n200_n840# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X709 fvf_1/Vbp bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X710 bbg_0/a_460_n780# fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X711 bbg_0/a_460_n780# bbg_0/a_460_n780# bbg_0/RES inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X712 fvf_1/VP fvf_1/Vbp bbg_0/a_460_n780# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X713 bbg_0/VBN bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X714 bbg_0/VBN bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X715 fvf_1/VP bbg_0/a_n200_n840# bbg_0/a_n200_n840# fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X716 inv_7/VN bbg_0/VBN fvf_1/Vbp inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X717 bbg_0/RES bbg_0/a_460_n780# bbg_0/a_460_n780# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X718 inv_7/VN bbg_0/VBN bbg_0/VBN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X719 fvf_1/VP bbg_0/a_n200_n840# fvf_1/Vbp fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X720 fvf_1/VP bbg_0/a_n200_n840# fvf_1/Vbp fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X721 inv_7/VN bbg_0/VBN bbg_0/VBN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X722 inv_7/VN bbg_0/a_460_n780# bbg_0/a_n200_n840# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X723 fvf_1/Vbp bbg_0/VBN inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X724 bbg_0/VBN fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X725 bbg_0/a_n200_n840# bbg_0/a_n200_n840# fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X726 fvf_0/Vin fvf_1/Vc fvf_0/Vdsg inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=1 ps=5 w=2 l=5
X727 fvf_0/Vin fvf_0/Vdsg inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=5
X728 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=1
X729 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=1
X730 fvf_0/Vdsg fvf_1/Vc fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0.5 ps=2.5 w=2 l=5
X731 fvf_0/Vdsg fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=1
X732 fvf_0/Vin fvf_1/Vc fvf_0/Vdsg inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=1 ps=5 w=2 l=5
X733 fvf_1/VP fvf_1/Vbp fvf_0/Vdsg fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1
X734 fvf_0/Vdsg fvf_1/Vc fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0.5 ps=2.5 w=2 l=5
X735 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=1
X736 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=1
X737 inv_7/VN fvf_0/Vdsg fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=5
X738 fvf_0/Vin fvf_0/Vdsg inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=5
X739 fvf_0/Vdsg fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=1
X740 fvf_1/VP fvf_1/Vbp fvf_0/Vdsg fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=1
X741 inv_7/VN fvf_0/Vdsg fvf_0/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=5
X742 fvf_1/Vin fvf_1/Vc Vcn inv_7/VN sky130_fd_pr__nfet_01v8 ad=9.25 pd=55 as=4 ps=20 w=2 l=5
X743 fvf_1/Vin Vcn inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=5
X744 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=1
X745 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=1
X746 Vcn fvf_1/Vc fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=5
X747 Vcn fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=2 pd=12 as=0 ps=0 w=1 l=1
X748 fvf_1/Vin fvf_1/Vc Vcn inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=5
X749 fvf_1/VP fvf_1/Vbp Vcn fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=1
X750 Vcn fvf_1/Vc fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=5
X751 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=1
X752 fvf_1/VP fvf_1/VP fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=1
X753 inv_7/VN Vcn fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=5
X754 fvf_1/Vin Vcn inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=5
X755 Vcn fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=1
X756 fvf_1/VP fvf_1/Vbp Vcn fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=1
X757 inv_7/VN Vcn fvf_1/Vin inv_7/VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=5
X758 inv_7/VN a_5360_22200# a_5360_22200# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=1
X759 inv_7/VN a_5360_22200# a_5360_22200# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=1
X760 inv_7/VP fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=3
X761 fvf_1/VP fvf_1/Vbp inv_7/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=3
X762 a_5360_22200# a_5360_22200# inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=1
X763 inv_7/VP inv_7/VP a_5360_22200# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=1
X764 a_5360_22200# inv_7/VP inv_7/VP inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=1
X765 inv_7/VP fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=3
X766 a_5360_22200# a_5360_22200# inv_7/VN inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=1
X767 fvf_1/VP fvf_1/Vbp inv_7/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.22 pd=1.9 as=0.22 ps=1.9 w=0.55 l=3
X768 dac_0/Iin fvf_1/Vbp fvf_1/VP fvf_1/VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=1
X769 inv_7/VP inv_7/VP a_5360_22200# inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=1
X770 a_5360_22200# inv_7/VP inv_7/VP inv_7/VN sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=1
